`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 22.05.2023 18:32:07
// Design Name: 
// Module Name: InstructionCache
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module InstructionCache(
    input clk,
    input [31:2] addr,
    output reg [31:0] data
    );
    
     // local variable
    wire addr_valid = (addr[31:14] == 18'h0);
    wire [11:0] dealt_addr = addr[13:2];
    // cache content
    reg [31:0] inst_cache [0:4095];
    
    
    always@(posedge clk)begin
        data <= addr_valid ? inst_cache[dealt_addr] : 32'h0;
    end
    
    initial begin
        data = 32'h0;
        inst_cache[       0] = 32'h00000013;
        inst_cache[       1] = 32'h00000093;
        inst_cache[       2] = 32'h00000113;
        inst_cache[       3] = 32'h00208f33;
        inst_cache[       4] = 32'h00000e93;
        inst_cache[       5] = 32'h00200193;
        inst_cache[       6] = 32'h01df0463;
        inst_cache[       7] = 32'h2ac0206f;
        inst_cache[       8] = 32'h00100093;
        inst_cache[       9] = 32'h00100113;
        inst_cache[      10] = 32'h00208f33;
        inst_cache[      11] = 32'h00200e93;
        inst_cache[      12] = 32'h00300193;
        inst_cache[      13] = 32'h01df0463;
        inst_cache[      14] = 32'h2900206f;
        inst_cache[      15] = 32'h00300093;
        inst_cache[      16] = 32'h00700113;
        inst_cache[      17] = 32'h00208f33;
        inst_cache[      18] = 32'h00a00e93;
        inst_cache[      19] = 32'h00400193;
        inst_cache[      20] = 32'h01df0463;
        inst_cache[      21] = 32'h2740206f;
        inst_cache[      22] = 32'h00000093;
        inst_cache[      23] = 32'hffff8137;
        inst_cache[      24] = 32'h00208f33;
        inst_cache[      25] = 32'hffff8eb7;
        inst_cache[      26] = 32'h00500193;
        inst_cache[      27] = 32'h01df0463;
        inst_cache[      28] = 32'h2580206f;
        inst_cache[      29] = 32'h800000b7;
        inst_cache[      30] = 32'h00000113;
        inst_cache[      31] = 32'h00208f33;
        inst_cache[      32] = 32'h80000eb7;
        inst_cache[      33] = 32'h00600193;
        inst_cache[      34] = 32'h01df0463;
        inst_cache[      35] = 32'h23c0206f;
        inst_cache[      36] = 32'h800000b7;
        inst_cache[      37] = 32'hffff8137;
        inst_cache[      38] = 32'h00208f33;
        inst_cache[      39] = 32'h7fff8eb7;
        inst_cache[      40] = 32'h00700193;
        inst_cache[      41] = 32'h01df0463;
        inst_cache[      42] = 32'h2200206f;
        inst_cache[      43] = 32'h00000093;
        inst_cache[      44] = 32'h00008137;
        inst_cache[      45] = 32'hfff10113;
        inst_cache[      46] = 32'h00208f33;
        inst_cache[      47] = 32'h00008eb7;
        inst_cache[      48] = 32'hfffe8e93;
        inst_cache[      49] = 32'h00800193;
        inst_cache[      50] = 32'h01df0463;
        inst_cache[      51] = 32'h1fc0206f;
        inst_cache[      52] = 32'h800000b7;
        inst_cache[      53] = 32'hfff08093;
        inst_cache[      54] = 32'h00000113;
        inst_cache[      55] = 32'h00208f33;
        inst_cache[      56] = 32'h80000eb7;
        inst_cache[      57] = 32'hfffe8e93;
        inst_cache[      58] = 32'h00900193;
        inst_cache[      59] = 32'h01df0463;
        inst_cache[      60] = 32'h1d80206f;
        inst_cache[      61] = 32'h800000b7;
        inst_cache[      62] = 32'hfff08093;
        inst_cache[      63] = 32'h00008137;
        inst_cache[      64] = 32'hfff10113;
        inst_cache[      65] = 32'h00208f33;
        inst_cache[      66] = 32'h80008eb7;
        inst_cache[      67] = 32'hffee8e93;
        inst_cache[      68] = 32'h00a00193;
        inst_cache[      69] = 32'h01df0463;
        inst_cache[      70] = 32'h1b00206f;
        inst_cache[      71] = 32'h800000b7;
        inst_cache[      72] = 32'h00008137;
        inst_cache[      73] = 32'hfff10113;
        inst_cache[      74] = 32'h00208f33;
        inst_cache[      75] = 32'h80008eb7;
        inst_cache[      76] = 32'hfffe8e93;
        inst_cache[      77] = 32'h00b00193;
        inst_cache[      78] = 32'h01df0463;
        inst_cache[      79] = 32'h18c0206f;
        inst_cache[      80] = 32'h800000b7;
        inst_cache[      81] = 32'hfff08093;
        inst_cache[      82] = 32'hffff8137;
        inst_cache[      83] = 32'h00208f33;
        inst_cache[      84] = 32'h7fff8eb7;
        inst_cache[      85] = 32'hfffe8e93;
        inst_cache[      86] = 32'h00c00193;
        inst_cache[      87] = 32'h01df0463;
        inst_cache[      88] = 32'h1680206f;
        inst_cache[      89] = 32'h00000093;
        inst_cache[      90] = 32'hfff00113;
        inst_cache[      91] = 32'h00208f33;
        inst_cache[      92] = 32'hfff00e93;
        inst_cache[      93] = 32'h00d00193;
        inst_cache[      94] = 32'h01df0463;
        inst_cache[      95] = 32'h14c0206f;
        inst_cache[      96] = 32'hfff00093;
        inst_cache[      97] = 32'h00100113;
        inst_cache[      98] = 32'h00208f33;
        inst_cache[      99] = 32'h00000e93;
        inst_cache[     100] = 32'h00e00193;
        inst_cache[     101] = 32'h01df0463;
        inst_cache[     102] = 32'h1300206f;
        inst_cache[     103] = 32'hfff00093;
        inst_cache[     104] = 32'hfff00113;
        inst_cache[     105] = 32'h00208f33;
        inst_cache[     106] = 32'hffe00e93;
        inst_cache[     107] = 32'h00f00193;
        inst_cache[     108] = 32'h01df0463;
        inst_cache[     109] = 32'h1140206f;
        inst_cache[     110] = 32'h00100093;
        inst_cache[     111] = 32'h80000137;
        inst_cache[     112] = 32'hfff10113;
        inst_cache[     113] = 32'h00208f33;
        inst_cache[     114] = 32'h80000eb7;
        inst_cache[     115] = 32'h01000193;
        inst_cache[     116] = 32'h01df0463;
        inst_cache[     117] = 32'h0f40206f;
        inst_cache[     118] = 32'h00d00093;
        inst_cache[     119] = 32'h00b00113;
        inst_cache[     120] = 32'h002080b3;
        inst_cache[     121] = 32'h01800e93;
        inst_cache[     122] = 32'h01100193;
        inst_cache[     123] = 32'h01d08463;
        inst_cache[     124] = 32'h0d80206f;
        inst_cache[     125] = 32'h00e00093;
        inst_cache[     126] = 32'h00b00113;
        inst_cache[     127] = 32'h00208133;
        inst_cache[     128] = 32'h01900e93;
        inst_cache[     129] = 32'h01200193;
        inst_cache[     130] = 32'h01d10463;
        inst_cache[     131] = 32'h0bc0206f;
        inst_cache[     132] = 32'h00d00093;
        inst_cache[     133] = 32'h001080b3;
        inst_cache[     134] = 32'h01a00e93;
        inst_cache[     135] = 32'h01300193;
        inst_cache[     136] = 32'h01d08463;
        inst_cache[     137] = 32'h0a40206f;
        inst_cache[     138] = 32'h00000213;
        inst_cache[     139] = 32'h00d00093;
        inst_cache[     140] = 32'h00b00113;
        inst_cache[     141] = 32'h00208f33;
        inst_cache[     142] = 32'h000f0313;
        inst_cache[     143] = 32'h00120213;
        inst_cache[     144] = 32'h00200293;
        inst_cache[     145] = 32'hfe5214e3;
        inst_cache[     146] = 32'h01800e93;
        inst_cache[     147] = 32'h01400193;
        inst_cache[     148] = 32'h01d30463;
        inst_cache[     149] = 32'h0740206f;
        inst_cache[     150] = 32'h00000213;
        inst_cache[     151] = 32'h00e00093;
        inst_cache[     152] = 32'h00b00113;
        inst_cache[     153] = 32'h00208f33;
        inst_cache[     154] = 32'h00000013;
        inst_cache[     155] = 32'h000f0313;
        inst_cache[     156] = 32'h00120213;
        inst_cache[     157] = 32'h00200293;
        inst_cache[     158] = 32'hfe5212e3;
        inst_cache[     159] = 32'h01900e93;
        inst_cache[     160] = 32'h01500193;
        inst_cache[     161] = 32'h01d30463;
        inst_cache[     162] = 32'h0400206f;
        inst_cache[     163] = 32'h00000213;
        inst_cache[     164] = 32'h00f00093;
        inst_cache[     165] = 32'h00b00113;
        inst_cache[     166] = 32'h00208f33;
        inst_cache[     167] = 32'h00000013;
        inst_cache[     168] = 32'h00000013;
        inst_cache[     169] = 32'h000f0313;
        inst_cache[     170] = 32'h00120213;
        inst_cache[     171] = 32'h00200293;
        inst_cache[     172] = 32'hfe5210e3;
        inst_cache[     173] = 32'h01a00e93;
        inst_cache[     174] = 32'h01600193;
        inst_cache[     175] = 32'h01d30463;
        inst_cache[     176] = 32'h0080206f;
        inst_cache[     177] = 32'h00000213;
        inst_cache[     178] = 32'h00d00093;
        inst_cache[     179] = 32'h00b00113;
        inst_cache[     180] = 32'h00208f33;
        inst_cache[     181] = 32'h00120213;
        inst_cache[     182] = 32'h00200293;
        inst_cache[     183] = 32'hfe5216e3;
        inst_cache[     184] = 32'h01800e93;
        inst_cache[     185] = 32'h01700193;
        inst_cache[     186] = 32'h01df0463;
        inst_cache[     187] = 32'h7dd0106f;
        inst_cache[     188] = 32'h00000213;
        inst_cache[     189] = 32'h00e00093;
        inst_cache[     190] = 32'h00b00113;
        inst_cache[     191] = 32'h00000013;
        inst_cache[     192] = 32'h00208f33;
        inst_cache[     193] = 32'h00120213;
        inst_cache[     194] = 32'h00200293;
        inst_cache[     195] = 32'hfe5214e3;
        inst_cache[     196] = 32'h01900e93;
        inst_cache[     197] = 32'h01800193;
        inst_cache[     198] = 32'h01df0463;
        inst_cache[     199] = 32'h7ad0106f;
        inst_cache[     200] = 32'h00000213;
        inst_cache[     201] = 32'h00f00093;
        inst_cache[     202] = 32'h00b00113;
        inst_cache[     203] = 32'h00000013;
        inst_cache[     204] = 32'h00000013;
        inst_cache[     205] = 32'h00208f33;
        inst_cache[     206] = 32'h00120213;
        inst_cache[     207] = 32'h00200293;
        inst_cache[     208] = 32'hfe5212e3;
        inst_cache[     209] = 32'h01a00e93;
        inst_cache[     210] = 32'h01900193;
        inst_cache[     211] = 32'h01df0463;
        inst_cache[     212] = 32'h7790106f;
        inst_cache[     213] = 32'h00000213;
        inst_cache[     214] = 32'h00d00093;
        inst_cache[     215] = 32'h00000013;
        inst_cache[     216] = 32'h00b00113;
        inst_cache[     217] = 32'h00208f33;
        inst_cache[     218] = 32'h00120213;
        inst_cache[     219] = 32'h00200293;
        inst_cache[     220] = 32'hfe5214e3;
        inst_cache[     221] = 32'h01800e93;
        inst_cache[     222] = 32'h01a00193;
        inst_cache[     223] = 32'h01df0463;
        inst_cache[     224] = 32'h7490106f;
        inst_cache[     225] = 32'h00000213;
        inst_cache[     226] = 32'h00e00093;
        inst_cache[     227] = 32'h00000013;
        inst_cache[     228] = 32'h00b00113;
        inst_cache[     229] = 32'h00000013;
        inst_cache[     230] = 32'h00208f33;
        inst_cache[     231] = 32'h00120213;
        inst_cache[     232] = 32'h00200293;
        inst_cache[     233] = 32'hfe5212e3;
        inst_cache[     234] = 32'h01900e93;
        inst_cache[     235] = 32'h01b00193;
        inst_cache[     236] = 32'h01df0463;
        inst_cache[     237] = 32'h7150106f;
        inst_cache[     238] = 32'h00000213;
        inst_cache[     239] = 32'h00f00093;
        inst_cache[     240] = 32'h00000013;
        inst_cache[     241] = 32'h00000013;
        inst_cache[     242] = 32'h00b00113;
        inst_cache[     243] = 32'h00208f33;
        inst_cache[     244] = 32'h00120213;
        inst_cache[     245] = 32'h00200293;
        inst_cache[     246] = 32'hfe5212e3;
        inst_cache[     247] = 32'h01a00e93;
        inst_cache[     248] = 32'h01c00193;
        inst_cache[     249] = 32'h01df0463;
        inst_cache[     250] = 32'h6e10106f;
        inst_cache[     251] = 32'h00000213;
        inst_cache[     252] = 32'h00b00113;
        inst_cache[     253] = 32'h00d00093;
        inst_cache[     254] = 32'h00208f33;
        inst_cache[     255] = 32'h00120213;
        inst_cache[     256] = 32'h00200293;
        inst_cache[     257] = 32'hfe5216e3;
        inst_cache[     258] = 32'h01800e93;
        inst_cache[     259] = 32'h01d00193;
        inst_cache[     260] = 32'h01df0463;
        inst_cache[     261] = 32'h6b50106f;
        inst_cache[     262] = 32'h00000213;
        inst_cache[     263] = 32'h00b00113;
        inst_cache[     264] = 32'h00e00093;
        inst_cache[     265] = 32'h00000013;
        inst_cache[     266] = 32'h00208f33;
        inst_cache[     267] = 32'h00120213;
        inst_cache[     268] = 32'h00200293;
        inst_cache[     269] = 32'hfe5214e3;
        inst_cache[     270] = 32'h01900e93;
        inst_cache[     271] = 32'h01e00193;
        inst_cache[     272] = 32'h01df0463;
        inst_cache[     273] = 32'h6850106f;
        inst_cache[     274] = 32'h00000213;
        inst_cache[     275] = 32'h00b00113;
        inst_cache[     276] = 32'h00f00093;
        inst_cache[     277] = 32'h00000013;
        inst_cache[     278] = 32'h00000013;
        inst_cache[     279] = 32'h00208f33;
        inst_cache[     280] = 32'h00120213;
        inst_cache[     281] = 32'h00200293;
        inst_cache[     282] = 32'hfe5212e3;
        inst_cache[     283] = 32'h01a00e93;
        inst_cache[     284] = 32'h01f00193;
        inst_cache[     285] = 32'h01df0463;
        inst_cache[     286] = 32'h6510106f;
        inst_cache[     287] = 32'h00000213;
        inst_cache[     288] = 32'h00b00113;
        inst_cache[     289] = 32'h00000013;
        inst_cache[     290] = 32'h00d00093;
        inst_cache[     291] = 32'h00208f33;
        inst_cache[     292] = 32'h00120213;
        inst_cache[     293] = 32'h00200293;
        inst_cache[     294] = 32'hfe5214e3;
        inst_cache[     295] = 32'h01800e93;
        inst_cache[     296] = 32'h02000193;
        inst_cache[     297] = 32'h01df0463;
        inst_cache[     298] = 32'h6210106f;
        inst_cache[     299] = 32'h00000213;
        inst_cache[     300] = 32'h00b00113;
        inst_cache[     301] = 32'h00000013;
        inst_cache[     302] = 32'h00e00093;
        inst_cache[     303] = 32'h00000013;
        inst_cache[     304] = 32'h00208f33;
        inst_cache[     305] = 32'h00120213;
        inst_cache[     306] = 32'h00200293;
        inst_cache[     307] = 32'hfe5212e3;
        inst_cache[     308] = 32'h01900e93;
        inst_cache[     309] = 32'h02100193;
        inst_cache[     310] = 32'h01df0463;
        inst_cache[     311] = 32'h5ed0106f;
        inst_cache[     312] = 32'h00000213;
        inst_cache[     313] = 32'h00b00113;
        inst_cache[     314] = 32'h00000013;
        inst_cache[     315] = 32'h00000013;
        inst_cache[     316] = 32'h00f00093;
        inst_cache[     317] = 32'h00208f33;
        inst_cache[     318] = 32'h00120213;
        inst_cache[     319] = 32'h00200293;
        inst_cache[     320] = 32'hfe5212e3;
        inst_cache[     321] = 32'h01a00e93;
        inst_cache[     322] = 32'h02200193;
        inst_cache[     323] = 32'h01df0463;
        inst_cache[     324] = 32'h5b90106f;
        inst_cache[     325] = 32'h00f00093;
        inst_cache[     326] = 32'h00100133;
        inst_cache[     327] = 32'h00f00e93;
        inst_cache[     328] = 32'h02300193;
        inst_cache[     329] = 32'h01d10463;
        inst_cache[     330] = 32'h5a10106f;
        inst_cache[     331] = 32'h02000093;
        inst_cache[     332] = 32'h00008133;
        inst_cache[     333] = 32'h02000e93;
        inst_cache[     334] = 32'h02400193;
        inst_cache[     335] = 32'h01d10463;
        inst_cache[     336] = 32'h5890106f;
        inst_cache[     337] = 32'h000000b3;
        inst_cache[     338] = 32'h00000e93;
        inst_cache[     339] = 32'h02500193;
        inst_cache[     340] = 32'h01d08463;
        inst_cache[     341] = 32'h5750106f;
        inst_cache[     342] = 32'h01000093;
        inst_cache[     343] = 32'h01e00113;
        inst_cache[     344] = 32'h00208033;
        inst_cache[     345] = 32'h00000e93;
        inst_cache[     346] = 32'h02600193;
        inst_cache[     347] = 32'h01d00463;
        inst_cache[     348] = 32'h5590106f;
        inst_cache[     349] = 32'h00000093;
        inst_cache[     350] = 32'h00008f13;
        inst_cache[     351] = 32'h00000e93;
        inst_cache[     352] = 32'h02700193;
        inst_cache[     353] = 32'h01df0463;
        inst_cache[     354] = 32'h5410106f;
        inst_cache[     355] = 32'h00100093;
        inst_cache[     356] = 32'h00108f13;
        inst_cache[     357] = 32'h00200e93;
        inst_cache[     358] = 32'h02800193;
        inst_cache[     359] = 32'h01df0463;
        inst_cache[     360] = 32'h5290106f;
        inst_cache[     361] = 32'h00300093;
        inst_cache[     362] = 32'h00708f13;
        inst_cache[     363] = 32'h00a00e93;
        inst_cache[     364] = 32'h02900193;
        inst_cache[     365] = 32'h01df0463;
        inst_cache[     366] = 32'h5110106f;
        inst_cache[     367] = 32'h00000093;
        inst_cache[     368] = 32'h80008f13;
        inst_cache[     369] = 32'h80000e93;
        inst_cache[     370] = 32'h02a00193;
        inst_cache[     371] = 32'h01df0463;
        inst_cache[     372] = 32'h4f90106f;
        inst_cache[     373] = 32'h800000b7;
        inst_cache[     374] = 32'h00008f13;
        inst_cache[     375] = 32'h80000eb7;
        inst_cache[     376] = 32'h02b00193;
        inst_cache[     377] = 32'h01df0463;
        inst_cache[     378] = 32'h4e10106f;
        inst_cache[     379] = 32'h800000b7;
        inst_cache[     380] = 32'h80008f13;
        inst_cache[     381] = 32'h80000eb7;
        inst_cache[     382] = 32'h800e8e93;
        inst_cache[     383] = 32'h02c00193;
        inst_cache[     384] = 32'h01df0463;
        inst_cache[     385] = 32'h4c50106f;
        inst_cache[     386] = 32'h00000093;
        inst_cache[     387] = 32'h7ff08f13;
        inst_cache[     388] = 32'h7ff00e93;
        inst_cache[     389] = 32'h02d00193;
        inst_cache[     390] = 32'h01df0463;
        inst_cache[     391] = 32'h4ad0106f;
        inst_cache[     392] = 32'h800000b7;
        inst_cache[     393] = 32'hfff08093;
        inst_cache[     394] = 32'h00008f13;
        inst_cache[     395] = 32'h80000eb7;
        inst_cache[     396] = 32'hfffe8e93;
        inst_cache[     397] = 32'h02e00193;
        inst_cache[     398] = 32'h01df0463;
        inst_cache[     399] = 32'h48d0106f;
        inst_cache[     400] = 32'h800000b7;
        inst_cache[     401] = 32'hfff08093;
        inst_cache[     402] = 32'h7ff08f13;
        inst_cache[     403] = 32'h80000eb7;
        inst_cache[     404] = 32'h7fee8e93;
        inst_cache[     405] = 32'h02f00193;
        inst_cache[     406] = 32'h01df0463;
        inst_cache[     407] = 32'h46d0106f;
        inst_cache[     408] = 32'h800000b7;
        inst_cache[     409] = 32'h7ff08f13;
        inst_cache[     410] = 32'h80000eb7;
        inst_cache[     411] = 32'h7ffe8e93;
        inst_cache[     412] = 32'h03000193;
        inst_cache[     413] = 32'h01df0463;
        inst_cache[     414] = 32'h4510106f;
        inst_cache[     415] = 32'h800000b7;
        inst_cache[     416] = 32'hfff08093;
        inst_cache[     417] = 32'h80008f13;
        inst_cache[     418] = 32'h7ffffeb7;
        inst_cache[     419] = 32'h7ffe8e93;
        inst_cache[     420] = 32'h03100193;
        inst_cache[     421] = 32'h01df0463;
        inst_cache[     422] = 32'h4310106f;
        inst_cache[     423] = 32'h00000093;
        inst_cache[     424] = 32'hfff08f13;
        inst_cache[     425] = 32'hfff00e93;
        inst_cache[     426] = 32'h03200193;
        inst_cache[     427] = 32'h01df0463;
        inst_cache[     428] = 32'h4190106f;
        inst_cache[     429] = 32'hfff00093;
        inst_cache[     430] = 32'h00108f13;
        inst_cache[     431] = 32'h00000e93;
        inst_cache[     432] = 32'h03300193;
        inst_cache[     433] = 32'h01df0463;
        inst_cache[     434] = 32'h4010106f;
        inst_cache[     435] = 32'hfff00093;
        inst_cache[     436] = 32'hfff08f13;
        inst_cache[     437] = 32'hffe00e93;
        inst_cache[     438] = 32'h03400193;
        inst_cache[     439] = 32'h01df0463;
        inst_cache[     440] = 32'h3e90106f;
        inst_cache[     441] = 32'h800000b7;
        inst_cache[     442] = 32'hfff08093;
        inst_cache[     443] = 32'h00108f13;
        inst_cache[     444] = 32'h80000eb7;
        inst_cache[     445] = 32'h03500193;
        inst_cache[     446] = 32'h01df0463;
        inst_cache[     447] = 32'h3cd0106f;
        inst_cache[     448] = 32'h00d00093;
        inst_cache[     449] = 32'h00b08093;
        inst_cache[     450] = 32'h01800e93;
        inst_cache[     451] = 32'h03600193;
        inst_cache[     452] = 32'h01d08463;
        inst_cache[     453] = 32'h3b50106f;
        inst_cache[     454] = 32'h00000213;
        inst_cache[     455] = 32'h00d00093;
        inst_cache[     456] = 32'h00b08f13;
        inst_cache[     457] = 32'h000f0313;
        inst_cache[     458] = 32'h00120213;
        inst_cache[     459] = 32'h00200293;
        inst_cache[     460] = 32'hfe5216e3;
        inst_cache[     461] = 32'h01800e93;
        inst_cache[     462] = 32'h03700193;
        inst_cache[     463] = 32'h01d30463;
        inst_cache[     464] = 32'h3890106f;
        inst_cache[     465] = 32'h00000213;
        inst_cache[     466] = 32'h00d00093;
        inst_cache[     467] = 32'h00a08f13;
        inst_cache[     468] = 32'h00000013;
        inst_cache[     469] = 32'h000f0313;
        inst_cache[     470] = 32'h00120213;
        inst_cache[     471] = 32'h00200293;
        inst_cache[     472] = 32'hfe5214e3;
        inst_cache[     473] = 32'h01700e93;
        inst_cache[     474] = 32'h03800193;
        inst_cache[     475] = 32'h01d30463;
        inst_cache[     476] = 32'h3590106f;
        inst_cache[     477] = 32'h00000213;
        inst_cache[     478] = 32'h00d00093;
        inst_cache[     479] = 32'h00908f13;
        inst_cache[     480] = 32'h00000013;
        inst_cache[     481] = 32'h00000013;
        inst_cache[     482] = 32'h000f0313;
        inst_cache[     483] = 32'h00120213;
        inst_cache[     484] = 32'h00200293;
        inst_cache[     485] = 32'hfe5212e3;
        inst_cache[     486] = 32'h01600e93;
        inst_cache[     487] = 32'h03900193;
        inst_cache[     488] = 32'h01d30463;
        inst_cache[     489] = 32'h3250106f;
        inst_cache[     490] = 32'h00000213;
        inst_cache[     491] = 32'h00d00093;
        inst_cache[     492] = 32'h00b08f13;
        inst_cache[     493] = 32'h00120213;
        inst_cache[     494] = 32'h00200293;
        inst_cache[     495] = 32'hfe5218e3;
        inst_cache[     496] = 32'h01800e93;
        inst_cache[     497] = 32'h03a00193;
        inst_cache[     498] = 32'h01df0463;
        inst_cache[     499] = 32'h2fd0106f;
        inst_cache[     500] = 32'h00000213;
        inst_cache[     501] = 32'h00d00093;
        inst_cache[     502] = 32'h00000013;
        inst_cache[     503] = 32'h00a08f13;
        inst_cache[     504] = 32'h00120213;
        inst_cache[     505] = 32'h00200293;
        inst_cache[     506] = 32'hfe5216e3;
        inst_cache[     507] = 32'h01700e93;
        inst_cache[     508] = 32'h03b00193;
        inst_cache[     509] = 32'h01df0463;
        inst_cache[     510] = 32'h2d10106f;
        inst_cache[     511] = 32'h00000213;
        inst_cache[     512] = 32'h00d00093;
        inst_cache[     513] = 32'h00000013;
        inst_cache[     514] = 32'h00000013;
        inst_cache[     515] = 32'h00908f13;
        inst_cache[     516] = 32'h00120213;
        inst_cache[     517] = 32'h00200293;
        inst_cache[     518] = 32'hfe5214e3;
        inst_cache[     519] = 32'h01600e93;
        inst_cache[     520] = 32'h03c00193;
        inst_cache[     521] = 32'h01df0463;
        inst_cache[     522] = 32'h2a10106f;
        inst_cache[     523] = 32'h02000093;
        inst_cache[     524] = 32'h02000e93;
        inst_cache[     525] = 32'h03d00193;
        inst_cache[     526] = 32'h01d08463;
        inst_cache[     527] = 32'h28d0106f;
        inst_cache[     528] = 32'h02100093;
        inst_cache[     529] = 32'h03208013;
        inst_cache[     530] = 32'h00000e93;
        inst_cache[     531] = 32'h03e00193;
        inst_cache[     532] = 32'h01d00463;
        inst_cache[     533] = 32'h2750106f;
        inst_cache[     534] = 32'hff0100b7;
        inst_cache[     535] = 32'hf0008093;
        inst_cache[     536] = 32'h0f0f1137;
        inst_cache[     537] = 32'hf0f10113;
        inst_cache[     538] = 32'h0020ff33;
        inst_cache[     539] = 32'h0f001eb7;
        inst_cache[     540] = 32'hf00e8e93;
        inst_cache[     541] = 32'h03f00193;
        inst_cache[     542] = 32'h01df0463;
        inst_cache[     543] = 32'h24d0106f;
        inst_cache[     544] = 32'h0ff010b7;
        inst_cache[     545] = 32'hff008093;
        inst_cache[     546] = 32'hf0f0f137;
        inst_cache[     547] = 32'h0f010113;
        inst_cache[     548] = 32'h0020ff33;
        inst_cache[     549] = 32'h00f00eb7;
        inst_cache[     550] = 32'h0f0e8e93;
        inst_cache[     551] = 32'h04000193;
        inst_cache[     552] = 32'h01df0463;
        inst_cache[     553] = 32'h2250106f;
        inst_cache[     554] = 32'h00ff00b7;
        inst_cache[     555] = 32'h0ff08093;
        inst_cache[     556] = 32'h0f0f1137;
        inst_cache[     557] = 32'hf0f10113;
        inst_cache[     558] = 32'h0020ff33;
        inst_cache[     559] = 32'h000f0eb7;
        inst_cache[     560] = 32'h00fe8e93;
        inst_cache[     561] = 32'h04100193;
        inst_cache[     562] = 32'h01df0463;
        inst_cache[     563] = 32'h1fd0106f;
        inst_cache[     564] = 32'hf00ff0b7;
        inst_cache[     565] = 32'h00f08093;
        inst_cache[     566] = 32'hf0f0f137;
        inst_cache[     567] = 32'h0f010113;
        inst_cache[     568] = 32'h0020ff33;
        inst_cache[     569] = 32'hf000feb7;
        inst_cache[     570] = 32'h04200193;
        inst_cache[     571] = 32'h01df0463;
        inst_cache[     572] = 32'h1d90106f;
        inst_cache[     573] = 32'hff0100b7;
        inst_cache[     574] = 32'hf0008093;
        inst_cache[     575] = 32'h0f0f1137;
        inst_cache[     576] = 32'hf0f10113;
        inst_cache[     577] = 32'h0020f0b3;
        inst_cache[     578] = 32'h0f001eb7;
        inst_cache[     579] = 32'hf00e8e93;
        inst_cache[     580] = 32'h04300193;
        inst_cache[     581] = 32'h01d08463;
        inst_cache[     582] = 32'h1b10106f;
        inst_cache[     583] = 32'h0ff010b7;
        inst_cache[     584] = 32'hff008093;
        inst_cache[     585] = 32'hf0f0f137;
        inst_cache[     586] = 32'h0f010113;
        inst_cache[     587] = 32'h0020f133;
        inst_cache[     588] = 32'h00f00eb7;
        inst_cache[     589] = 32'h0f0e8e93;
        inst_cache[     590] = 32'h04400193;
        inst_cache[     591] = 32'h01d10463;
        inst_cache[     592] = 32'h1890106f;
        inst_cache[     593] = 32'hff0100b7;
        inst_cache[     594] = 32'hf0008093;
        inst_cache[     595] = 32'h0010f0b3;
        inst_cache[     596] = 32'hff010eb7;
        inst_cache[     597] = 32'hf00e8e93;
        inst_cache[     598] = 32'h04500193;
        inst_cache[     599] = 32'h01d08463;
        inst_cache[     600] = 32'h1690106f;
        inst_cache[     601] = 32'h00000213;
        inst_cache[     602] = 32'hff0100b7;
        inst_cache[     603] = 32'hf0008093;
        inst_cache[     604] = 32'h0f0f1137;
        inst_cache[     605] = 32'hf0f10113;
        inst_cache[     606] = 32'h0020ff33;
        inst_cache[     607] = 32'h000f0313;
        inst_cache[     608] = 32'h00120213;
        inst_cache[     609] = 32'h00200293;
        inst_cache[     610] = 32'hfe5210e3;
        inst_cache[     611] = 32'h0f001eb7;
        inst_cache[     612] = 32'hf00e8e93;
        inst_cache[     613] = 32'h04600193;
        inst_cache[     614] = 32'h01d30463;
        inst_cache[     615] = 32'h12d0106f;
        inst_cache[     616] = 32'h00000213;
        inst_cache[     617] = 32'h0ff010b7;
        inst_cache[     618] = 32'hff008093;
        inst_cache[     619] = 32'hf0f0f137;
        inst_cache[     620] = 32'h0f010113;
        inst_cache[     621] = 32'h0020ff33;
        inst_cache[     622] = 32'h00000013;
        inst_cache[     623] = 32'h000f0313;
        inst_cache[     624] = 32'h00120213;
        inst_cache[     625] = 32'h00200293;
        inst_cache[     626] = 32'hfc521ee3;
        inst_cache[     627] = 32'h00f00eb7;
        inst_cache[     628] = 32'h0f0e8e93;
        inst_cache[     629] = 32'h04700193;
        inst_cache[     630] = 32'h01d30463;
        inst_cache[     631] = 32'h0ed0106f;
        inst_cache[     632] = 32'h00000213;
        inst_cache[     633] = 32'h00ff00b7;
        inst_cache[     634] = 32'h0ff08093;
        inst_cache[     635] = 32'h0f0f1137;
        inst_cache[     636] = 32'hf0f10113;
        inst_cache[     637] = 32'h0020ff33;
        inst_cache[     638] = 32'h00000013;
        inst_cache[     639] = 32'h00000013;
        inst_cache[     640] = 32'h000f0313;
        inst_cache[     641] = 32'h00120213;
        inst_cache[     642] = 32'h00200293;
        inst_cache[     643] = 32'hfc521ce3;
        inst_cache[     644] = 32'h000f0eb7;
        inst_cache[     645] = 32'h00fe8e93;
        inst_cache[     646] = 32'h04800193;
        inst_cache[     647] = 32'h01d30463;
        inst_cache[     648] = 32'h0a90106f;
        inst_cache[     649] = 32'h00000213;
        inst_cache[     650] = 32'hff0100b7;
        inst_cache[     651] = 32'hf0008093;
        inst_cache[     652] = 32'h0f0f1137;
        inst_cache[     653] = 32'hf0f10113;
        inst_cache[     654] = 32'h0020ff33;
        inst_cache[     655] = 32'h00120213;
        inst_cache[     656] = 32'h00200293;
        inst_cache[     657] = 32'hfe5212e3;
        inst_cache[     658] = 32'h0f001eb7;
        inst_cache[     659] = 32'hf00e8e93;
        inst_cache[     660] = 32'h04900193;
        inst_cache[     661] = 32'h01df0463;
        inst_cache[     662] = 32'h0710106f;
        inst_cache[     663] = 32'h00000213;
        inst_cache[     664] = 32'h0ff010b7;
        inst_cache[     665] = 32'hff008093;
        inst_cache[     666] = 32'hf0f0f137;
        inst_cache[     667] = 32'h0f010113;
        inst_cache[     668] = 32'h00000013;
        inst_cache[     669] = 32'h0020ff33;
        inst_cache[     670] = 32'h00120213;
        inst_cache[     671] = 32'h00200293;
        inst_cache[     672] = 32'hfe5210e3;
        inst_cache[     673] = 32'h00f00eb7;
        inst_cache[     674] = 32'h0f0e8e93;
        inst_cache[     675] = 32'h04a00193;
        inst_cache[     676] = 32'h01df0463;
        inst_cache[     677] = 32'h0350106f;
        inst_cache[     678] = 32'h00000213;
        inst_cache[     679] = 32'h00ff00b7;
        inst_cache[     680] = 32'h0ff08093;
        inst_cache[     681] = 32'h0f0f1137;
        inst_cache[     682] = 32'hf0f10113;
        inst_cache[     683] = 32'h00000013;
        inst_cache[     684] = 32'h00000013;
        inst_cache[     685] = 32'h0020ff33;
        inst_cache[     686] = 32'h00120213;
        inst_cache[     687] = 32'h00200293;
        inst_cache[     688] = 32'hfc521ee3;
        inst_cache[     689] = 32'h000f0eb7;
        inst_cache[     690] = 32'h00fe8e93;
        inst_cache[     691] = 32'h04b00193;
        inst_cache[     692] = 32'h01df0463;
        inst_cache[     693] = 32'h7f40106f;
        inst_cache[     694] = 32'h00000213;
        inst_cache[     695] = 32'hff0100b7;
        inst_cache[     696] = 32'hf0008093;
        inst_cache[     697] = 32'h00000013;
        inst_cache[     698] = 32'h0f0f1137;
        inst_cache[     699] = 32'hf0f10113;
        inst_cache[     700] = 32'h0020ff33;
        inst_cache[     701] = 32'h00120213;
        inst_cache[     702] = 32'h00200293;
        inst_cache[     703] = 32'hfe5210e3;
        inst_cache[     704] = 32'h0f001eb7;
        inst_cache[     705] = 32'hf00e8e93;
        inst_cache[     706] = 32'h04c00193;
        inst_cache[     707] = 32'h01df0463;
        inst_cache[     708] = 32'h7b80106f;
        inst_cache[     709] = 32'h00000213;
        inst_cache[     710] = 32'h0ff010b7;
        inst_cache[     711] = 32'hff008093;
        inst_cache[     712] = 32'h00000013;
        inst_cache[     713] = 32'hf0f0f137;
        inst_cache[     714] = 32'h0f010113;
        inst_cache[     715] = 32'h00000013;
        inst_cache[     716] = 32'h0020ff33;
        inst_cache[     717] = 32'h00120213;
        inst_cache[     718] = 32'h00200293;
        inst_cache[     719] = 32'hfc521ee3;
        inst_cache[     720] = 32'h00f00eb7;
        inst_cache[     721] = 32'h0f0e8e93;
        inst_cache[     722] = 32'h04d00193;
        inst_cache[     723] = 32'h01df0463;
        inst_cache[     724] = 32'h7780106f;
        inst_cache[     725] = 32'h00000213;
        inst_cache[     726] = 32'h00ff00b7;
        inst_cache[     727] = 32'h0ff08093;
        inst_cache[     728] = 32'h00000013;
        inst_cache[     729] = 32'h00000013;
        inst_cache[     730] = 32'h0f0f1137;
        inst_cache[     731] = 32'hf0f10113;
        inst_cache[     732] = 32'h0020ff33;
        inst_cache[     733] = 32'h00120213;
        inst_cache[     734] = 32'h00200293;
        inst_cache[     735] = 32'hfc521ee3;
        inst_cache[     736] = 32'h000f0eb7;
        inst_cache[     737] = 32'h00fe8e93;
        inst_cache[     738] = 32'h04e00193;
        inst_cache[     739] = 32'h01df0463;
        inst_cache[     740] = 32'h7380106f;
        inst_cache[     741] = 32'h00000213;
        inst_cache[     742] = 32'h0f0f1137;
        inst_cache[     743] = 32'hf0f10113;
        inst_cache[     744] = 32'hff0100b7;
        inst_cache[     745] = 32'hf0008093;
        inst_cache[     746] = 32'h0020ff33;
        inst_cache[     747] = 32'h00120213;
        inst_cache[     748] = 32'h00200293;
        inst_cache[     749] = 32'hfe5212e3;
        inst_cache[     750] = 32'h0f001eb7;
        inst_cache[     751] = 32'hf00e8e93;
        inst_cache[     752] = 32'h04f00193;
        inst_cache[     753] = 32'h01df0463;
        inst_cache[     754] = 32'h7000106f;
        inst_cache[     755] = 32'h00000213;
        inst_cache[     756] = 32'hf0f0f137;
        inst_cache[     757] = 32'h0f010113;
        inst_cache[     758] = 32'h0ff010b7;
        inst_cache[     759] = 32'hff008093;
        inst_cache[     760] = 32'h00000013;
        inst_cache[     761] = 32'h0020ff33;
        inst_cache[     762] = 32'h00120213;
        inst_cache[     763] = 32'h00200293;
        inst_cache[     764] = 32'hfe5210e3;
        inst_cache[     765] = 32'h00f00eb7;
        inst_cache[     766] = 32'h0f0e8e93;
        inst_cache[     767] = 32'h05000193;
        inst_cache[     768] = 32'h01df0463;
        inst_cache[     769] = 32'h6c40106f;
        inst_cache[     770] = 32'h00000213;
        inst_cache[     771] = 32'h0f0f1137;
        inst_cache[     772] = 32'hf0f10113;
        inst_cache[     773] = 32'h00ff00b7;
        inst_cache[     774] = 32'h0ff08093;
        inst_cache[     775] = 32'h00000013;
        inst_cache[     776] = 32'h00000013;
        inst_cache[     777] = 32'h0020ff33;
        inst_cache[     778] = 32'h00120213;
        inst_cache[     779] = 32'h00200293;
        inst_cache[     780] = 32'hfc521ee3;
        inst_cache[     781] = 32'h000f0eb7;
        inst_cache[     782] = 32'h00fe8e93;
        inst_cache[     783] = 32'h05100193;
        inst_cache[     784] = 32'h01df0463;
        inst_cache[     785] = 32'h6840106f;
        inst_cache[     786] = 32'h00000213;
        inst_cache[     787] = 32'h0f0f1137;
        inst_cache[     788] = 32'hf0f10113;
        inst_cache[     789] = 32'h00000013;
        inst_cache[     790] = 32'hff0100b7;
        inst_cache[     791] = 32'hf0008093;
        inst_cache[     792] = 32'h0020ff33;
        inst_cache[     793] = 32'h00120213;
        inst_cache[     794] = 32'h00200293;
        inst_cache[     795] = 32'hfe5210e3;
        inst_cache[     796] = 32'h0f001eb7;
        inst_cache[     797] = 32'hf00e8e93;
        inst_cache[     798] = 32'h05200193;
        inst_cache[     799] = 32'h01df0463;
        inst_cache[     800] = 32'h6480106f;
        inst_cache[     801] = 32'h00000213;
        inst_cache[     802] = 32'hf0f0f137;
        inst_cache[     803] = 32'h0f010113;
        inst_cache[     804] = 32'h00000013;
        inst_cache[     805] = 32'h0ff010b7;
        inst_cache[     806] = 32'hff008093;
        inst_cache[     807] = 32'h00000013;
        inst_cache[     808] = 32'h0020ff33;
        inst_cache[     809] = 32'h00120213;
        inst_cache[     810] = 32'h00200293;
        inst_cache[     811] = 32'hfc521ee3;
        inst_cache[     812] = 32'h00f00eb7;
        inst_cache[     813] = 32'h0f0e8e93;
        inst_cache[     814] = 32'h05300193;
        inst_cache[     815] = 32'h01df0463;
        inst_cache[     816] = 32'h6080106f;
        inst_cache[     817] = 32'h00000213;
        inst_cache[     818] = 32'h0f0f1137;
        inst_cache[     819] = 32'hf0f10113;
        inst_cache[     820] = 32'h00000013;
        inst_cache[     821] = 32'h00000013;
        inst_cache[     822] = 32'h00ff00b7;
        inst_cache[     823] = 32'h0ff08093;
        inst_cache[     824] = 32'h0020ff33;
        inst_cache[     825] = 32'h00120213;
        inst_cache[     826] = 32'h00200293;
        inst_cache[     827] = 32'hfc521ee3;
        inst_cache[     828] = 32'h000f0eb7;
        inst_cache[     829] = 32'h00fe8e93;
        inst_cache[     830] = 32'h05400193;
        inst_cache[     831] = 32'h01df0463;
        inst_cache[     832] = 32'h5c80106f;
        inst_cache[     833] = 32'hff0100b7;
        inst_cache[     834] = 32'hf0008093;
        inst_cache[     835] = 32'h00107133;
        inst_cache[     836] = 32'h00000e93;
        inst_cache[     837] = 32'h05500193;
        inst_cache[     838] = 32'h01d10463;
        inst_cache[     839] = 32'h5ac0106f;
        inst_cache[     840] = 32'h00ff00b7;
        inst_cache[     841] = 32'h0ff08093;
        inst_cache[     842] = 32'h0000f133;
        inst_cache[     843] = 32'h00000e93;
        inst_cache[     844] = 32'h05600193;
        inst_cache[     845] = 32'h01d10463;
        inst_cache[     846] = 32'h5900106f;
        inst_cache[     847] = 32'h000070b3;
        inst_cache[     848] = 32'h00000e93;
        inst_cache[     849] = 32'h05700193;
        inst_cache[     850] = 32'h01d08463;
        inst_cache[     851] = 32'h57c0106f;
        inst_cache[     852] = 32'h111110b7;
        inst_cache[     853] = 32'h11108093;
        inst_cache[     854] = 32'h22222137;
        inst_cache[     855] = 32'h22210113;
        inst_cache[     856] = 32'h0020f033;
        inst_cache[     857] = 32'h00000e93;
        inst_cache[     858] = 32'h05800193;
        inst_cache[     859] = 32'h01d00463;
        inst_cache[     860] = 32'h5580106f;
        inst_cache[     861] = 32'hff0100b7;
        inst_cache[     862] = 32'hf0008093;
        inst_cache[     863] = 32'hf0f0ff13;
        inst_cache[     864] = 32'hff010eb7;
        inst_cache[     865] = 32'hf00e8e93;
        inst_cache[     866] = 32'h05900193;
        inst_cache[     867] = 32'h01df0463;
        inst_cache[     868] = 32'h5380106f;
        inst_cache[     869] = 32'h0ff010b7;
        inst_cache[     870] = 32'hff008093;
        inst_cache[     871] = 32'h0f00ff13;
        inst_cache[     872] = 32'h0f000e93;
        inst_cache[     873] = 32'h05a00193;
        inst_cache[     874] = 32'h01df0463;
        inst_cache[     875] = 32'h51c0106f;
        inst_cache[     876] = 32'h00ff00b7;
        inst_cache[     877] = 32'h0ff08093;
        inst_cache[     878] = 32'h70f0ff13;
        inst_cache[     879] = 32'h00f00e93;
        inst_cache[     880] = 32'h05b00193;
        inst_cache[     881] = 32'h01df0463;
        inst_cache[     882] = 32'h5000106f;
        inst_cache[     883] = 32'hf00ff0b7;
        inst_cache[     884] = 32'h00f08093;
        inst_cache[     885] = 32'h0f00ff13;
        inst_cache[     886] = 32'h00000e93;
        inst_cache[     887] = 32'h05c00193;
        inst_cache[     888] = 32'h01df0463;
        inst_cache[     889] = 32'h4e40106f;
        inst_cache[     890] = 32'hff0100b7;
        inst_cache[     891] = 32'hf0008093;
        inst_cache[     892] = 32'h0f00f093;
        inst_cache[     893] = 32'h00000e93;
        inst_cache[     894] = 32'h05d00193;
        inst_cache[     895] = 32'h01d08463;
        inst_cache[     896] = 32'h4c80106f;
        inst_cache[     897] = 32'h00000213;
        inst_cache[     898] = 32'h0ff010b7;
        inst_cache[     899] = 32'hff008093;
        inst_cache[     900] = 32'h70f0ff13;
        inst_cache[     901] = 32'h000f0313;
        inst_cache[     902] = 32'h00120213;
        inst_cache[     903] = 32'h00200293;
        inst_cache[     904] = 32'hfe5214e3;
        inst_cache[     905] = 32'h70000e93;
        inst_cache[     906] = 32'h05e00193;
        inst_cache[     907] = 32'h01d30463;
        inst_cache[     908] = 32'h4980106f;
        inst_cache[     909] = 32'h00000213;
        inst_cache[     910] = 32'h00ff00b7;
        inst_cache[     911] = 32'h0ff08093;
        inst_cache[     912] = 32'h0f00ff13;
        inst_cache[     913] = 32'h00000013;
        inst_cache[     914] = 32'h000f0313;
        inst_cache[     915] = 32'h00120213;
        inst_cache[     916] = 32'h00200293;
        inst_cache[     917] = 32'hfe5212e3;
        inst_cache[     918] = 32'h0f000e93;
        inst_cache[     919] = 32'h05f00193;
        inst_cache[     920] = 32'h01d30463;
        inst_cache[     921] = 32'h4640106f;
        inst_cache[     922] = 32'h00000213;
        inst_cache[     923] = 32'hf00ff0b7;
        inst_cache[     924] = 32'h00f08093;
        inst_cache[     925] = 32'hf0f0ff13;
        inst_cache[     926] = 32'h00000013;
        inst_cache[     927] = 32'h00000013;
        inst_cache[     928] = 32'h000f0313;
        inst_cache[     929] = 32'h00120213;
        inst_cache[     930] = 32'h00200293;
        inst_cache[     931] = 32'hfe5210e3;
        inst_cache[     932] = 32'hf00ffeb7;
        inst_cache[     933] = 32'h00fe8e93;
        inst_cache[     934] = 32'h06000193;
        inst_cache[     935] = 32'h01d30463;
        inst_cache[     936] = 32'h4280106f;
        inst_cache[     937] = 32'h00000213;
        inst_cache[     938] = 32'h0ff010b7;
        inst_cache[     939] = 32'hff008093;
        inst_cache[     940] = 32'h70f0ff13;
        inst_cache[     941] = 32'h00120213;
        inst_cache[     942] = 32'h00200293;
        inst_cache[     943] = 32'hfe5216e3;
        inst_cache[     944] = 32'h70000e93;
        inst_cache[     945] = 32'h06100193;
        inst_cache[     946] = 32'h01df0463;
        inst_cache[     947] = 32'h3fc0106f;
        inst_cache[     948] = 32'h00000213;
        inst_cache[     949] = 32'h00ff00b7;
        inst_cache[     950] = 32'h0ff08093;
        inst_cache[     951] = 32'h00000013;
        inst_cache[     952] = 32'h0f00ff13;
        inst_cache[     953] = 32'h00120213;
        inst_cache[     954] = 32'h00200293;
        inst_cache[     955] = 32'hfe5214e3;
        inst_cache[     956] = 32'h0f000e93;
        inst_cache[     957] = 32'h06200193;
        inst_cache[     958] = 32'h01df0463;
        inst_cache[     959] = 32'h3cc0106f;
        inst_cache[     960] = 32'h00000213;
        inst_cache[     961] = 32'hf00ff0b7;
        inst_cache[     962] = 32'h00f08093;
        inst_cache[     963] = 32'h00000013;
        inst_cache[     964] = 32'h00000013;
        inst_cache[     965] = 32'h70f0ff13;
        inst_cache[     966] = 32'h00120213;
        inst_cache[     967] = 32'h00200293;
        inst_cache[     968] = 32'hfe5212e3;
        inst_cache[     969] = 32'h00f00e93;
        inst_cache[     970] = 32'h06300193;
        inst_cache[     971] = 32'h01df0463;
        inst_cache[     972] = 32'h3980106f;
        inst_cache[     973] = 32'h0f007093;
        inst_cache[     974] = 32'h00000e93;
        inst_cache[     975] = 32'h06400193;
        inst_cache[     976] = 32'h01d08463;
        inst_cache[     977] = 32'h3840106f;
        inst_cache[     978] = 32'h00ff00b7;
        inst_cache[     979] = 32'h0ff08093;
        inst_cache[     980] = 32'h70f0f013;
        inst_cache[     981] = 32'h00000e93;
        inst_cache[     982] = 32'h06500193;
        inst_cache[     983] = 32'h01d00463;
        inst_cache[     984] = 32'h3680106f;
        inst_cache[     985] = 32'h00000013;
        inst_cache[     986] = 32'h00002517;
        inst_cache[     987] = 32'h71c50513;
        inst_cache[     988] = 32'h004005ef;
        inst_cache[     989] = 32'h40b50533;
        inst_cache[     990] = 32'h00002eb7;
        inst_cache[     991] = 32'h710e8e93;
        inst_cache[     992] = 32'h06600193;
        inst_cache[     993] = 32'h01d50463;
        inst_cache[     994] = 32'h3400106f;
        inst_cache[     995] = 32'h00000013;
        inst_cache[     996] = 32'hffffe517;
        inst_cache[     997] = 32'h8fc50513;
        inst_cache[     998] = 32'h004005ef;
        inst_cache[     999] = 32'h40b50533;
        inst_cache[    1000] = 32'hffffeeb7;
        inst_cache[    1001] = 32'h8f0e8e93;
        inst_cache[    1002] = 32'h06700193;
        inst_cache[    1003] = 32'h01d50463;
        inst_cache[    1004] = 32'h3180106f;
        inst_cache[    1005] = 32'h06800193;
        inst_cache[    1006] = 32'h00000093;
        inst_cache[    1007] = 32'h00000113;
        inst_cache[    1008] = 32'h00208863;
        inst_cache[    1009] = 32'h00300463;
        inst_cache[    1010] = 32'h3000106f;
        inst_cache[    1011] = 32'h00301863;
        inst_cache[    1012] = 32'hfe208ee3;
        inst_cache[    1013] = 32'h00300463;
        inst_cache[    1014] = 32'h2f00106f;
        inst_cache[    1015] = 32'h06900193;
        inst_cache[    1016] = 32'h00100093;
        inst_cache[    1017] = 32'h00100113;
        inst_cache[    1018] = 32'h00208863;
        inst_cache[    1019] = 32'h00300463;
        inst_cache[    1020] = 32'h2d80106f;
        inst_cache[    1021] = 32'h00301863;
        inst_cache[    1022] = 32'hfe208ee3;
        inst_cache[    1023] = 32'h00300463;
        inst_cache[    1024] = 32'h2c80106f;
        inst_cache[    1025] = 32'h06a00193;
        inst_cache[    1026] = 32'hfff00093;
        inst_cache[    1027] = 32'hfff00113;
        inst_cache[    1028] = 32'h00208863;
        inst_cache[    1029] = 32'h00300463;
        inst_cache[    1030] = 32'h2b00106f;
        inst_cache[    1031] = 32'h00301863;
        inst_cache[    1032] = 32'hfe208ee3;
        inst_cache[    1033] = 32'h00300463;
        inst_cache[    1034] = 32'h2a00106f;
        inst_cache[    1035] = 32'h06b00193;
        inst_cache[    1036] = 32'h00000093;
        inst_cache[    1037] = 32'h00100113;
        inst_cache[    1038] = 32'h00208463;
        inst_cache[    1039] = 32'h00301663;
        inst_cache[    1040] = 32'h00300463;
        inst_cache[    1041] = 32'h2840106f;
        inst_cache[    1042] = 32'hfe208ce3;
        inst_cache[    1043] = 32'h06c00193;
        inst_cache[    1044] = 32'h00100093;
        inst_cache[    1045] = 32'h00000113;
        inst_cache[    1046] = 32'h00208463;
        inst_cache[    1047] = 32'h00301663;
        inst_cache[    1048] = 32'h00300463;
        inst_cache[    1049] = 32'h2640106f;
        inst_cache[    1050] = 32'hfe208ce3;
        inst_cache[    1051] = 32'h06d00193;
        inst_cache[    1052] = 32'hfff00093;
        inst_cache[    1053] = 32'h00100113;
        inst_cache[    1054] = 32'h00208463;
        inst_cache[    1055] = 32'h00301663;
        inst_cache[    1056] = 32'h00300463;
        inst_cache[    1057] = 32'h2440106f;
        inst_cache[    1058] = 32'hfe208ce3;
        inst_cache[    1059] = 32'h06e00193;
        inst_cache[    1060] = 32'h00100093;
        inst_cache[    1061] = 32'hfff00113;
        inst_cache[    1062] = 32'h00208463;
        inst_cache[    1063] = 32'h00301663;
        inst_cache[    1064] = 32'h00300463;
        inst_cache[    1065] = 32'h2240106f;
        inst_cache[    1066] = 32'hfe208ce3;
        inst_cache[    1067] = 32'h06f00193;
        inst_cache[    1068] = 32'h00000213;
        inst_cache[    1069] = 32'h00000093;
        inst_cache[    1070] = 32'hfff00113;
        inst_cache[    1071] = 32'h00209463;
        inst_cache[    1072] = 32'h2080106f;
        inst_cache[    1073] = 32'h00120213;
        inst_cache[    1074] = 32'h00200293;
        inst_cache[    1075] = 32'hfe5214e3;
        inst_cache[    1076] = 32'h07000193;
        inst_cache[    1077] = 32'h00000213;
        inst_cache[    1078] = 32'h00000093;
        inst_cache[    1079] = 32'hfff00113;
        inst_cache[    1080] = 32'h00000013;
        inst_cache[    1081] = 32'h00209463;
        inst_cache[    1082] = 32'h1e00106f;
        inst_cache[    1083] = 32'h00120213;
        inst_cache[    1084] = 32'h00200293;
        inst_cache[    1085] = 32'hfe5212e3;
        inst_cache[    1086] = 32'h07100193;
        inst_cache[    1087] = 32'h00000213;
        inst_cache[    1088] = 32'h00000093;
        inst_cache[    1089] = 32'hfff00113;
        inst_cache[    1090] = 32'h00000013;
        inst_cache[    1091] = 32'h00000013;
        inst_cache[    1092] = 32'h00209463;
        inst_cache[    1093] = 32'h1b40106f;
        inst_cache[    1094] = 32'h00120213;
        inst_cache[    1095] = 32'h00200293;
        inst_cache[    1096] = 32'hfe5210e3;
        inst_cache[    1097] = 32'h07200193;
        inst_cache[    1098] = 32'h00000213;
        inst_cache[    1099] = 32'h00000093;
        inst_cache[    1100] = 32'h00000013;
        inst_cache[    1101] = 32'hfff00113;
        inst_cache[    1102] = 32'h00209463;
        inst_cache[    1103] = 32'h18c0106f;
        inst_cache[    1104] = 32'h00120213;
        inst_cache[    1105] = 32'h00200293;
        inst_cache[    1106] = 32'hfe5212e3;
        inst_cache[    1107] = 32'h07300193;
        inst_cache[    1108] = 32'h00000213;
        inst_cache[    1109] = 32'h00000093;
        inst_cache[    1110] = 32'h00000013;
        inst_cache[    1111] = 32'hfff00113;
        inst_cache[    1112] = 32'h00000013;
        inst_cache[    1113] = 32'h00209463;
        inst_cache[    1114] = 32'h1600106f;
        inst_cache[    1115] = 32'h00120213;
        inst_cache[    1116] = 32'h00200293;
        inst_cache[    1117] = 32'hfe5210e3;
        inst_cache[    1118] = 32'h07400193;
        inst_cache[    1119] = 32'h00000213;
        inst_cache[    1120] = 32'h00000093;
        inst_cache[    1121] = 32'h00000013;
        inst_cache[    1122] = 32'h00000013;
        inst_cache[    1123] = 32'hfff00113;
        inst_cache[    1124] = 32'h00209463;
        inst_cache[    1125] = 32'h1340106f;
        inst_cache[    1126] = 32'h00120213;
        inst_cache[    1127] = 32'h00200293;
        inst_cache[    1128] = 32'hfe5210e3;
        inst_cache[    1129] = 32'h07500193;
        inst_cache[    1130] = 32'h00000213;
        inst_cache[    1131] = 32'h00000093;
        inst_cache[    1132] = 32'hfff00113;
        inst_cache[    1133] = 32'h00209463;
        inst_cache[    1134] = 32'h1100106f;
        inst_cache[    1135] = 32'h00120213;
        inst_cache[    1136] = 32'h00200293;
        inst_cache[    1137] = 32'hfe5214e3;
        inst_cache[    1138] = 32'h07600193;
        inst_cache[    1139] = 32'h00000213;
        inst_cache[    1140] = 32'h00000093;
        inst_cache[    1141] = 32'hfff00113;
        inst_cache[    1142] = 32'h00000013;
        inst_cache[    1143] = 32'h00209463;
        inst_cache[    1144] = 32'h0e80106f;
        inst_cache[    1145] = 32'h00120213;
        inst_cache[    1146] = 32'h00200293;
        inst_cache[    1147] = 32'hfe5212e3;
        inst_cache[    1148] = 32'h07700193;
        inst_cache[    1149] = 32'h00000213;
        inst_cache[    1150] = 32'h00000093;
        inst_cache[    1151] = 32'hfff00113;
        inst_cache[    1152] = 32'h00000013;
        inst_cache[    1153] = 32'h00000013;
        inst_cache[    1154] = 32'h00209463;
        inst_cache[    1155] = 32'h0bc0106f;
        inst_cache[    1156] = 32'h00120213;
        inst_cache[    1157] = 32'h00200293;
        inst_cache[    1158] = 32'hfe5210e3;
        inst_cache[    1159] = 32'h07800193;
        inst_cache[    1160] = 32'h00000213;
        inst_cache[    1161] = 32'h00000093;
        inst_cache[    1162] = 32'h00000013;
        inst_cache[    1163] = 32'hfff00113;
        inst_cache[    1164] = 32'h00209463;
        inst_cache[    1165] = 32'h0940106f;
        inst_cache[    1166] = 32'h00120213;
        inst_cache[    1167] = 32'h00200293;
        inst_cache[    1168] = 32'hfe5212e3;
        inst_cache[    1169] = 32'h07900193;
        inst_cache[    1170] = 32'h00000213;
        inst_cache[    1171] = 32'h00000093;
        inst_cache[    1172] = 32'h00000013;
        inst_cache[    1173] = 32'hfff00113;
        inst_cache[    1174] = 32'h00000013;
        inst_cache[    1175] = 32'h00209463;
        inst_cache[    1176] = 32'h0680106f;
        inst_cache[    1177] = 32'h00120213;
        inst_cache[    1178] = 32'h00200293;
        inst_cache[    1179] = 32'hfe5210e3;
        inst_cache[    1180] = 32'h07a00193;
        inst_cache[    1181] = 32'h00000213;
        inst_cache[    1182] = 32'h00000093;
        inst_cache[    1183] = 32'h00000013;
        inst_cache[    1184] = 32'h00000013;
        inst_cache[    1185] = 32'hfff00113;
        inst_cache[    1186] = 32'h00209463;
        inst_cache[    1187] = 32'h03c0106f;
        inst_cache[    1188] = 32'h00120213;
        inst_cache[    1189] = 32'h00200293;
        inst_cache[    1190] = 32'hfe5210e3;
        inst_cache[    1191] = 32'h00100093;
        inst_cache[    1192] = 32'h00000a63;
        inst_cache[    1193] = 32'h00108093;
        inst_cache[    1194] = 32'h00108093;
        inst_cache[    1195] = 32'h00108093;
        inst_cache[    1196] = 32'h00108093;
        inst_cache[    1197] = 32'h00108093;
        inst_cache[    1198] = 32'h00108093;
        inst_cache[    1199] = 32'h00300e93;
        inst_cache[    1200] = 32'h07b00193;
        inst_cache[    1201] = 32'h01d08463;
        inst_cache[    1202] = 32'h0000106f;
        inst_cache[    1203] = 32'h07c00193;
        inst_cache[    1204] = 32'h00000093;
        inst_cache[    1205] = 32'h00000113;
        inst_cache[    1206] = 32'h0020d663;
        inst_cache[    1207] = 32'h7e3016e3;
        inst_cache[    1208] = 32'h00301663;
        inst_cache[    1209] = 32'hfe20dee3;
        inst_cache[    1210] = 32'h7e3010e3;
        inst_cache[    1211] = 32'h07d00193;
        inst_cache[    1212] = 32'h00100093;
        inst_cache[    1213] = 32'h00100113;
        inst_cache[    1214] = 32'h0020d663;
        inst_cache[    1215] = 32'h7c3016e3;
        inst_cache[    1216] = 32'h00301663;
        inst_cache[    1217] = 32'hfe20dee3;
        inst_cache[    1218] = 32'h7c3010e3;
        inst_cache[    1219] = 32'h07e00193;
        inst_cache[    1220] = 32'hfff00093;
        inst_cache[    1221] = 32'hfff00113;
        inst_cache[    1222] = 32'h0020d663;
        inst_cache[    1223] = 32'h7a3016e3;
        inst_cache[    1224] = 32'h00301663;
        inst_cache[    1225] = 32'hfe20dee3;
        inst_cache[    1226] = 32'h7a3010e3;
        inst_cache[    1227] = 32'h07f00193;
        inst_cache[    1228] = 32'h00100093;
        inst_cache[    1229] = 32'h00000113;
        inst_cache[    1230] = 32'h0020d663;
        inst_cache[    1231] = 32'h783016e3;
        inst_cache[    1232] = 32'h00301663;
        inst_cache[    1233] = 32'hfe20dee3;
        inst_cache[    1234] = 32'h783010e3;
        inst_cache[    1235] = 32'h08000193;
        inst_cache[    1236] = 32'h00100093;
        inst_cache[    1237] = 32'hfff00113;
        inst_cache[    1238] = 32'h0020d663;
        inst_cache[    1239] = 32'h763016e3;
        inst_cache[    1240] = 32'h00301663;
        inst_cache[    1241] = 32'hfe20dee3;
        inst_cache[    1242] = 32'h763010e3;
        inst_cache[    1243] = 32'h08100193;
        inst_cache[    1244] = 32'hfff00093;
        inst_cache[    1245] = 32'hffe00113;
        inst_cache[    1246] = 32'h0020d663;
        inst_cache[    1247] = 32'h743016e3;
        inst_cache[    1248] = 32'h00301663;
        inst_cache[    1249] = 32'hfe20dee3;
        inst_cache[    1250] = 32'h743010e3;
        inst_cache[    1251] = 32'h08200193;
        inst_cache[    1252] = 32'h00000093;
        inst_cache[    1253] = 32'h00100113;
        inst_cache[    1254] = 32'h0020d463;
        inst_cache[    1255] = 32'h00301463;
        inst_cache[    1256] = 32'h723014e3;
        inst_cache[    1257] = 32'hfe20dee3;
        inst_cache[    1258] = 32'h08300193;
        inst_cache[    1259] = 32'hfff00093;
        inst_cache[    1260] = 32'h00100113;
        inst_cache[    1261] = 32'h0020d463;
        inst_cache[    1262] = 32'h00301463;
        inst_cache[    1263] = 32'h703016e3;
        inst_cache[    1264] = 32'hfe20dee3;
        inst_cache[    1265] = 32'h08400193;
        inst_cache[    1266] = 32'hffe00093;
        inst_cache[    1267] = 32'hfff00113;
        inst_cache[    1268] = 32'h0020d463;
        inst_cache[    1269] = 32'h00301463;
        inst_cache[    1270] = 32'h6e3018e3;
        inst_cache[    1271] = 32'hfe20dee3;
        inst_cache[    1272] = 32'h08500193;
        inst_cache[    1273] = 32'hffe00093;
        inst_cache[    1274] = 32'h00100113;
        inst_cache[    1275] = 32'h0020d463;
        inst_cache[    1276] = 32'h00301463;
        inst_cache[    1277] = 32'h6c301ae3;
        inst_cache[    1278] = 32'hfe20dee3;
        inst_cache[    1279] = 32'h08600193;
        inst_cache[    1280] = 32'h00000213;
        inst_cache[    1281] = 32'hfff00093;
        inst_cache[    1282] = 32'h00000113;
        inst_cache[    1283] = 32'h6a20dee3;
        inst_cache[    1284] = 32'h00120213;
        inst_cache[    1285] = 32'h00200293;
        inst_cache[    1286] = 32'hfe5216e3;
        inst_cache[    1287] = 32'h08700193;
        inst_cache[    1288] = 32'h00000213;
        inst_cache[    1289] = 32'hfff00093;
        inst_cache[    1290] = 32'h00000113;
        inst_cache[    1291] = 32'h00000013;
        inst_cache[    1292] = 32'h6820dce3;
        inst_cache[    1293] = 32'h00120213;
        inst_cache[    1294] = 32'h00200293;
        inst_cache[    1295] = 32'hfe5214e3;
        inst_cache[    1296] = 32'h08800193;
        inst_cache[    1297] = 32'h00000213;
        inst_cache[    1298] = 32'hfff00093;
        inst_cache[    1299] = 32'h00000113;
        inst_cache[    1300] = 32'h00000013;
        inst_cache[    1301] = 32'h00000013;
        inst_cache[    1302] = 32'h6620d8e3;
        inst_cache[    1303] = 32'h00120213;
        inst_cache[    1304] = 32'h00200293;
        inst_cache[    1305] = 32'hfe5212e3;
        inst_cache[    1306] = 32'h08900193;
        inst_cache[    1307] = 32'h00000213;
        inst_cache[    1308] = 32'hfff00093;
        inst_cache[    1309] = 32'h00000013;
        inst_cache[    1310] = 32'h00000113;
        inst_cache[    1311] = 32'h6420d6e3;
        inst_cache[    1312] = 32'h00120213;
        inst_cache[    1313] = 32'h00200293;
        inst_cache[    1314] = 32'hfe5214e3;
        inst_cache[    1315] = 32'h08a00193;
        inst_cache[    1316] = 32'h00000213;
        inst_cache[    1317] = 32'hfff00093;
        inst_cache[    1318] = 32'h00000013;
        inst_cache[    1319] = 32'h00000113;
        inst_cache[    1320] = 32'h00000013;
        inst_cache[    1321] = 32'h6220d2e3;
        inst_cache[    1322] = 32'h00120213;
        inst_cache[    1323] = 32'h00200293;
        inst_cache[    1324] = 32'hfe5212e3;
        inst_cache[    1325] = 32'h08b00193;
        inst_cache[    1326] = 32'h00000213;
        inst_cache[    1327] = 32'hfff00093;
        inst_cache[    1328] = 32'h00000013;
        inst_cache[    1329] = 32'h00000013;
        inst_cache[    1330] = 32'h00000113;
        inst_cache[    1331] = 32'h5e20dee3;
        inst_cache[    1332] = 32'h00120213;
        inst_cache[    1333] = 32'h00200293;
        inst_cache[    1334] = 32'hfe5212e3;
        inst_cache[    1335] = 32'h08c00193;
        inst_cache[    1336] = 32'h00000213;
        inst_cache[    1337] = 32'hfff00093;
        inst_cache[    1338] = 32'h00000113;
        inst_cache[    1339] = 32'h5c20dee3;
        inst_cache[    1340] = 32'h00120213;
        inst_cache[    1341] = 32'h00200293;
        inst_cache[    1342] = 32'hfe5216e3;
        inst_cache[    1343] = 32'h08d00193;
        inst_cache[    1344] = 32'h00000213;
        inst_cache[    1345] = 32'hfff00093;
        inst_cache[    1346] = 32'h00000113;
        inst_cache[    1347] = 32'h00000013;
        inst_cache[    1348] = 32'h5a20dce3;
        inst_cache[    1349] = 32'h00120213;
        inst_cache[    1350] = 32'h00200293;
        inst_cache[    1351] = 32'hfe5214e3;
        inst_cache[    1352] = 32'h08e00193;
        inst_cache[    1353] = 32'h00000213;
        inst_cache[    1354] = 32'hfff00093;
        inst_cache[    1355] = 32'h00000113;
        inst_cache[    1356] = 32'h00000013;
        inst_cache[    1357] = 32'h00000013;
        inst_cache[    1358] = 32'h5820d8e3;
        inst_cache[    1359] = 32'h00120213;
        inst_cache[    1360] = 32'h00200293;
        inst_cache[    1361] = 32'hfe5212e3;
        inst_cache[    1362] = 32'h08f00193;
        inst_cache[    1363] = 32'h00000213;
        inst_cache[    1364] = 32'hfff00093;
        inst_cache[    1365] = 32'h00000013;
        inst_cache[    1366] = 32'h00000113;
        inst_cache[    1367] = 32'h5620d6e3;
        inst_cache[    1368] = 32'h00120213;
        inst_cache[    1369] = 32'h00200293;
        inst_cache[    1370] = 32'hfe5214e3;
        inst_cache[    1371] = 32'h09000193;
        inst_cache[    1372] = 32'h00000213;
        inst_cache[    1373] = 32'hfff00093;
        inst_cache[    1374] = 32'h00000013;
        inst_cache[    1375] = 32'h00000113;
        inst_cache[    1376] = 32'h00000013;
        inst_cache[    1377] = 32'h5420d2e3;
        inst_cache[    1378] = 32'h00120213;
        inst_cache[    1379] = 32'h00200293;
        inst_cache[    1380] = 32'hfe5212e3;
        inst_cache[    1381] = 32'h09100193;
        inst_cache[    1382] = 32'h00000213;
        inst_cache[    1383] = 32'hfff00093;
        inst_cache[    1384] = 32'h00000013;
        inst_cache[    1385] = 32'h00000013;
        inst_cache[    1386] = 32'h00000113;
        inst_cache[    1387] = 32'h5020dee3;
        inst_cache[    1388] = 32'h00120213;
        inst_cache[    1389] = 32'h00200293;
        inst_cache[    1390] = 32'hfe5212e3;
        inst_cache[    1391] = 32'h00100093;
        inst_cache[    1392] = 32'h0000da63;
        inst_cache[    1393] = 32'h00108093;
        inst_cache[    1394] = 32'h00108093;
        inst_cache[    1395] = 32'h00108093;
        inst_cache[    1396] = 32'h00108093;
        inst_cache[    1397] = 32'h00108093;
        inst_cache[    1398] = 32'h00108093;
        inst_cache[    1399] = 32'h00300e93;
        inst_cache[    1400] = 32'h09200193;
        inst_cache[    1401] = 32'h4fd092e3;
        inst_cache[    1402] = 32'h09300193;
        inst_cache[    1403] = 32'h00000093;
        inst_cache[    1404] = 32'h00000113;
        inst_cache[    1405] = 32'h0020f663;
        inst_cache[    1406] = 32'h4c3018e3;
        inst_cache[    1407] = 32'h00301663;
        inst_cache[    1408] = 32'hfe20fee3;
        inst_cache[    1409] = 32'h4c3012e3;
        inst_cache[    1410] = 32'h09400193;
        inst_cache[    1411] = 32'h00100093;
        inst_cache[    1412] = 32'h00100113;
        inst_cache[    1413] = 32'h0020f663;
        inst_cache[    1414] = 32'h4a3018e3;
        inst_cache[    1415] = 32'h00301663;
        inst_cache[    1416] = 32'hfe20fee3;
        inst_cache[    1417] = 32'h4a3012e3;
        inst_cache[    1418] = 32'h09500193;
        inst_cache[    1419] = 32'hfff00093;
        inst_cache[    1420] = 32'hfff00113;
        inst_cache[    1421] = 32'h0020f663;
        inst_cache[    1422] = 32'h483018e3;
        inst_cache[    1423] = 32'h00301663;
        inst_cache[    1424] = 32'hfe20fee3;
        inst_cache[    1425] = 32'h483012e3;
        inst_cache[    1426] = 32'h09600193;
        inst_cache[    1427] = 32'h00100093;
        inst_cache[    1428] = 32'h00000113;
        inst_cache[    1429] = 32'h0020f663;
        inst_cache[    1430] = 32'h463018e3;
        inst_cache[    1431] = 32'h00301663;
        inst_cache[    1432] = 32'hfe20fee3;
        inst_cache[    1433] = 32'h463012e3;
        inst_cache[    1434] = 32'h09700193;
        inst_cache[    1435] = 32'hfff00093;
        inst_cache[    1436] = 32'hffe00113;
        inst_cache[    1437] = 32'h0020f663;
        inst_cache[    1438] = 32'h443018e3;
        inst_cache[    1439] = 32'h00301663;
        inst_cache[    1440] = 32'hfe20fee3;
        inst_cache[    1441] = 32'h443012e3;
        inst_cache[    1442] = 32'h09800193;
        inst_cache[    1443] = 32'hfff00093;
        inst_cache[    1444] = 32'h00000113;
        inst_cache[    1445] = 32'h0020f663;
        inst_cache[    1446] = 32'h423018e3;
        inst_cache[    1447] = 32'h00301663;
        inst_cache[    1448] = 32'hfe20fee3;
        inst_cache[    1449] = 32'h423012e3;
        inst_cache[    1450] = 32'h09900193;
        inst_cache[    1451] = 32'h00000093;
        inst_cache[    1452] = 32'h00100113;
        inst_cache[    1453] = 32'h0020f463;
        inst_cache[    1454] = 32'h00301463;
        inst_cache[    1455] = 32'h403016e3;
        inst_cache[    1456] = 32'hfe20fee3;
        inst_cache[    1457] = 32'h09a00193;
        inst_cache[    1458] = 32'hffe00093;
        inst_cache[    1459] = 32'hfff00113;
        inst_cache[    1460] = 32'h0020f463;
        inst_cache[    1461] = 32'h00301463;
        inst_cache[    1462] = 32'h3e3018e3;
        inst_cache[    1463] = 32'hfe20fee3;
        inst_cache[    1464] = 32'h09b00193;
        inst_cache[    1465] = 32'h00000093;
        inst_cache[    1466] = 32'hfff00113;
        inst_cache[    1467] = 32'h0020f463;
        inst_cache[    1468] = 32'h00301463;
        inst_cache[    1469] = 32'h3c301ae3;
        inst_cache[    1470] = 32'hfe20fee3;
        inst_cache[    1471] = 32'h09c00193;
        inst_cache[    1472] = 32'h800000b7;
        inst_cache[    1473] = 32'hfff08093;
        inst_cache[    1474] = 32'h80000137;
        inst_cache[    1475] = 32'h0020f463;
        inst_cache[    1476] = 32'h00301463;
        inst_cache[    1477] = 32'h3a301ae3;
        inst_cache[    1478] = 32'hfe20fee3;
        inst_cache[    1479] = 32'h09d00193;
        inst_cache[    1480] = 32'h00000213;
        inst_cache[    1481] = 32'hf00000b7;
        inst_cache[    1482] = 32'hfff08093;
        inst_cache[    1483] = 32'hf0000137;
        inst_cache[    1484] = 32'h3820fce3;
        inst_cache[    1485] = 32'h00120213;
        inst_cache[    1486] = 32'h00200293;
        inst_cache[    1487] = 32'hfe5214e3;
        inst_cache[    1488] = 32'h09e00193;
        inst_cache[    1489] = 32'h00000213;
        inst_cache[    1490] = 32'hf00000b7;
        inst_cache[    1491] = 32'hfff08093;
        inst_cache[    1492] = 32'hf0000137;
        inst_cache[    1493] = 32'h00000013;
        inst_cache[    1494] = 32'h3620f8e3;
        inst_cache[    1495] = 32'h00120213;
        inst_cache[    1496] = 32'h00200293;
        inst_cache[    1497] = 32'hfe5212e3;
        inst_cache[    1498] = 32'h09f00193;
        inst_cache[    1499] = 32'h00000213;
        inst_cache[    1500] = 32'hf00000b7;
        inst_cache[    1501] = 32'hfff08093;
        inst_cache[    1502] = 32'hf0000137;
        inst_cache[    1503] = 32'h00000013;
        inst_cache[    1504] = 32'h00000013;
        inst_cache[    1505] = 32'h3420f2e3;
        inst_cache[    1506] = 32'h00120213;
        inst_cache[    1507] = 32'h00200293;
        inst_cache[    1508] = 32'hfe5210e3;
        inst_cache[    1509] = 32'h0a000193;
        inst_cache[    1510] = 32'h00000213;
        inst_cache[    1511] = 32'hf00000b7;
        inst_cache[    1512] = 32'hfff08093;
        inst_cache[    1513] = 32'h00000013;
        inst_cache[    1514] = 32'hf0000137;
        inst_cache[    1515] = 32'h3020fee3;
        inst_cache[    1516] = 32'h00120213;
        inst_cache[    1517] = 32'h00200293;
        inst_cache[    1518] = 32'hfe5212e3;
        inst_cache[    1519] = 32'h0a100193;
        inst_cache[    1520] = 32'h00000213;
        inst_cache[    1521] = 32'hf00000b7;
        inst_cache[    1522] = 32'hfff08093;
        inst_cache[    1523] = 32'h00000013;
        inst_cache[    1524] = 32'hf0000137;
        inst_cache[    1525] = 32'h00000013;
        inst_cache[    1526] = 32'h2e20f8e3;
        inst_cache[    1527] = 32'h00120213;
        inst_cache[    1528] = 32'h00200293;
        inst_cache[    1529] = 32'hfe5210e3;
        inst_cache[    1530] = 32'h0a200193;
        inst_cache[    1531] = 32'h00000213;
        inst_cache[    1532] = 32'hf00000b7;
        inst_cache[    1533] = 32'hfff08093;
        inst_cache[    1534] = 32'h00000013;
        inst_cache[    1535] = 32'h00000013;
        inst_cache[    1536] = 32'hf0000137;
        inst_cache[    1537] = 32'h2c20f2e3;
        inst_cache[    1538] = 32'h00120213;
        inst_cache[    1539] = 32'h00200293;
        inst_cache[    1540] = 32'hfe5210e3;
        inst_cache[    1541] = 32'h0a300193;
        inst_cache[    1542] = 32'h00000213;
        inst_cache[    1543] = 32'hf00000b7;
        inst_cache[    1544] = 32'hfff08093;
        inst_cache[    1545] = 32'hf0000137;
        inst_cache[    1546] = 32'h2a20f0e3;
        inst_cache[    1547] = 32'h00120213;
        inst_cache[    1548] = 32'h00200293;
        inst_cache[    1549] = 32'hfe5214e3;
        inst_cache[    1550] = 32'h0a400193;
        inst_cache[    1551] = 32'h00000213;
        inst_cache[    1552] = 32'hf00000b7;
        inst_cache[    1553] = 32'hfff08093;
        inst_cache[    1554] = 32'hf0000137;
        inst_cache[    1555] = 32'h00000013;
        inst_cache[    1556] = 32'h2620fce3;
        inst_cache[    1557] = 32'h00120213;
        inst_cache[    1558] = 32'h00200293;
        inst_cache[    1559] = 32'hfe5212e3;
        inst_cache[    1560] = 32'h0a500193;
        inst_cache[    1561] = 32'h00000213;
        inst_cache[    1562] = 32'hf00000b7;
        inst_cache[    1563] = 32'hfff08093;
        inst_cache[    1564] = 32'hf0000137;
        inst_cache[    1565] = 32'h00000013;
        inst_cache[    1566] = 32'h00000013;
        inst_cache[    1567] = 32'h2420f6e3;
        inst_cache[    1568] = 32'h00120213;
        inst_cache[    1569] = 32'h00200293;
        inst_cache[    1570] = 32'hfe5210e3;
        inst_cache[    1571] = 32'h0a600193;
        inst_cache[    1572] = 32'h00000213;
        inst_cache[    1573] = 32'hf00000b7;
        inst_cache[    1574] = 32'hfff08093;
        inst_cache[    1575] = 32'h00000013;
        inst_cache[    1576] = 32'hf0000137;
        inst_cache[    1577] = 32'h2220f2e3;
        inst_cache[    1578] = 32'h00120213;
        inst_cache[    1579] = 32'h00200293;
        inst_cache[    1580] = 32'hfe5212e3;
        inst_cache[    1581] = 32'h0a700193;
        inst_cache[    1582] = 32'h00000213;
        inst_cache[    1583] = 32'hf00000b7;
        inst_cache[    1584] = 32'hfff08093;
        inst_cache[    1585] = 32'h00000013;
        inst_cache[    1586] = 32'hf0000137;
        inst_cache[    1587] = 32'h00000013;
        inst_cache[    1588] = 32'h1e20fce3;
        inst_cache[    1589] = 32'h00120213;
        inst_cache[    1590] = 32'h00200293;
        inst_cache[    1591] = 32'hfe5210e3;
        inst_cache[    1592] = 32'h0a800193;
        inst_cache[    1593] = 32'h00000213;
        inst_cache[    1594] = 32'hf00000b7;
        inst_cache[    1595] = 32'hfff08093;
        inst_cache[    1596] = 32'h00000013;
        inst_cache[    1597] = 32'h00000013;
        inst_cache[    1598] = 32'hf0000137;
        inst_cache[    1599] = 32'h1c20f6e3;
        inst_cache[    1600] = 32'h00120213;
        inst_cache[    1601] = 32'h00200293;
        inst_cache[    1602] = 32'hfe5210e3;
        inst_cache[    1603] = 32'h00100093;
        inst_cache[    1604] = 32'h0000fa63;
        inst_cache[    1605] = 32'h00108093;
        inst_cache[    1606] = 32'h00108093;
        inst_cache[    1607] = 32'h00108093;
        inst_cache[    1608] = 32'h00108093;
        inst_cache[    1609] = 32'h00108093;
        inst_cache[    1610] = 32'h00108093;
        inst_cache[    1611] = 32'h00300e93;
        inst_cache[    1612] = 32'h0a900193;
        inst_cache[    1613] = 32'h19d09ae3;
        inst_cache[    1614] = 32'h0aa00193;
        inst_cache[    1615] = 32'h00000093;
        inst_cache[    1616] = 32'h00100113;
        inst_cache[    1617] = 32'h0020c663;
        inst_cache[    1618] = 32'h183010e3;
        inst_cache[    1619] = 32'h00301663;
        inst_cache[    1620] = 32'hfe20cee3;
        inst_cache[    1621] = 32'h16301ae3;
        inst_cache[    1622] = 32'h0ab00193;
        inst_cache[    1623] = 32'hfff00093;
        inst_cache[    1624] = 32'h00100113;
        inst_cache[    1625] = 32'h0020c663;
        inst_cache[    1626] = 32'h163010e3;
        inst_cache[    1627] = 32'h00301663;
        inst_cache[    1628] = 32'hfe20cee3;
        inst_cache[    1629] = 32'h14301ae3;
        inst_cache[    1630] = 32'h0ac00193;
        inst_cache[    1631] = 32'hffe00093;
        inst_cache[    1632] = 32'hfff00113;
        inst_cache[    1633] = 32'h0020c663;
        inst_cache[    1634] = 32'h143010e3;
        inst_cache[    1635] = 32'h00301663;
        inst_cache[    1636] = 32'hfe20cee3;
        inst_cache[    1637] = 32'h12301ae3;
        inst_cache[    1638] = 32'h0ad00193;
        inst_cache[    1639] = 32'h00100093;
        inst_cache[    1640] = 32'h00000113;
        inst_cache[    1641] = 32'h0020c463;
        inst_cache[    1642] = 32'h00301463;
        inst_cache[    1643] = 32'h10301ee3;
        inst_cache[    1644] = 32'hfe20cee3;
        inst_cache[    1645] = 32'h0ae00193;
        inst_cache[    1646] = 32'h00100093;
        inst_cache[    1647] = 32'hfff00113;
        inst_cache[    1648] = 32'h0020c463;
        inst_cache[    1649] = 32'h00301463;
        inst_cache[    1650] = 32'h103010e3;
        inst_cache[    1651] = 32'hfe20cee3;
        inst_cache[    1652] = 32'h0af00193;
        inst_cache[    1653] = 32'hfff00093;
        inst_cache[    1654] = 32'hffe00113;
        inst_cache[    1655] = 32'h0020c463;
        inst_cache[    1656] = 32'h00301463;
        inst_cache[    1657] = 32'h0e3012e3;
        inst_cache[    1658] = 32'hfe20cee3;
        inst_cache[    1659] = 32'h0b000193;
        inst_cache[    1660] = 32'h00100093;
        inst_cache[    1661] = 32'hffe00113;
        inst_cache[    1662] = 32'h0020c463;
        inst_cache[    1663] = 32'h00301463;
        inst_cache[    1664] = 32'h0c3014e3;
        inst_cache[    1665] = 32'hfe20cee3;
        inst_cache[    1666] = 32'h0b100193;
        inst_cache[    1667] = 32'h00000213;
        inst_cache[    1668] = 32'h00000093;
        inst_cache[    1669] = 32'hfff00113;
        inst_cache[    1670] = 32'h0a20c8e3;
        inst_cache[    1671] = 32'h00120213;
        inst_cache[    1672] = 32'h00200293;
        inst_cache[    1673] = 32'hfe5216e3;
        inst_cache[    1674] = 32'h0b200193;
        inst_cache[    1675] = 32'h00000213;
        inst_cache[    1676] = 32'h00000093;
        inst_cache[    1677] = 32'hfff00113;
        inst_cache[    1678] = 32'h00000013;
        inst_cache[    1679] = 32'h0820c6e3;
        inst_cache[    1680] = 32'h00120213;
        inst_cache[    1681] = 32'h00200293;
        inst_cache[    1682] = 32'hfe5214e3;
        inst_cache[    1683] = 32'h0b300193;
        inst_cache[    1684] = 32'h00000213;
        inst_cache[    1685] = 32'h00000093;
        inst_cache[    1686] = 32'hfff00113;
        inst_cache[    1687] = 32'h00000013;
        inst_cache[    1688] = 32'h00000013;
        inst_cache[    1689] = 32'h0620c2e3;
        inst_cache[    1690] = 32'h00120213;
        inst_cache[    1691] = 32'h00200293;
        inst_cache[    1692] = 32'hfe5212e3;
        inst_cache[    1693] = 32'h0b400193;
        inst_cache[    1694] = 32'h00000213;
        inst_cache[    1695] = 32'h00000093;
        inst_cache[    1696] = 32'h00000013;
        inst_cache[    1697] = 32'hfff00113;
        inst_cache[    1698] = 32'h0420c0e3;
        inst_cache[    1699] = 32'h00120213;
        inst_cache[    1700] = 32'h00200293;
        inst_cache[    1701] = 32'hfe5214e3;
        inst_cache[    1702] = 32'h0b500193;
        inst_cache[    1703] = 32'h00000213;
        inst_cache[    1704] = 32'h00000093;
        inst_cache[    1705] = 32'h00000013;
        inst_cache[    1706] = 32'hfff00113;
        inst_cache[    1707] = 32'h00000013;
        inst_cache[    1708] = 32'h0020cce3;
        inst_cache[    1709] = 32'h00120213;
        inst_cache[    1710] = 32'h00200293;
        inst_cache[    1711] = 32'hfe5212e3;
        inst_cache[    1712] = 32'h0b600193;
        inst_cache[    1713] = 32'h00000213;
        inst_cache[    1714] = 32'h00000093;
        inst_cache[    1715] = 32'h00000013;
        inst_cache[    1716] = 32'h00000013;
        inst_cache[    1717] = 32'hfff00113;
        inst_cache[    1718] = 32'h7e20c863;
        inst_cache[    1719] = 32'h00120213;
        inst_cache[    1720] = 32'h00200293;
        inst_cache[    1721] = 32'hfe5212e3;
        inst_cache[    1722] = 32'h0b700193;
        inst_cache[    1723] = 32'h00000213;
        inst_cache[    1724] = 32'h00000093;
        inst_cache[    1725] = 32'hfff00113;
        inst_cache[    1726] = 32'h7c20c863;
        inst_cache[    1727] = 32'h00120213;
        inst_cache[    1728] = 32'h00200293;
        inst_cache[    1729] = 32'hfe5216e3;
        inst_cache[    1730] = 32'h0b800193;
        inst_cache[    1731] = 32'h00000213;
        inst_cache[    1732] = 32'h00000093;
        inst_cache[    1733] = 32'hfff00113;
        inst_cache[    1734] = 32'h00000013;
        inst_cache[    1735] = 32'h7a20c663;
        inst_cache[    1736] = 32'h00120213;
        inst_cache[    1737] = 32'h00200293;
        inst_cache[    1738] = 32'hfe5214e3;
        inst_cache[    1739] = 32'h0b900193;
        inst_cache[    1740] = 32'h00000213;
        inst_cache[    1741] = 32'h00000093;
        inst_cache[    1742] = 32'hfff00113;
        inst_cache[    1743] = 32'h00000013;
        inst_cache[    1744] = 32'h00000013;
        inst_cache[    1745] = 32'h7820c263;
        inst_cache[    1746] = 32'h00120213;
        inst_cache[    1747] = 32'h00200293;
        inst_cache[    1748] = 32'hfe5212e3;
        inst_cache[    1749] = 32'h0ba00193;
        inst_cache[    1750] = 32'h00000213;
        inst_cache[    1751] = 32'h00000093;
        inst_cache[    1752] = 32'h00000013;
        inst_cache[    1753] = 32'hfff00113;
        inst_cache[    1754] = 32'h7620c063;
        inst_cache[    1755] = 32'h00120213;
        inst_cache[    1756] = 32'h00200293;
        inst_cache[    1757] = 32'hfe5214e3;
        inst_cache[    1758] = 32'h0bb00193;
        inst_cache[    1759] = 32'h00000213;
        inst_cache[    1760] = 32'h00000093;
        inst_cache[    1761] = 32'h00000013;
        inst_cache[    1762] = 32'hfff00113;
        inst_cache[    1763] = 32'h00000013;
        inst_cache[    1764] = 32'h7220cc63;
        inst_cache[    1765] = 32'h00120213;
        inst_cache[    1766] = 32'h00200293;
        inst_cache[    1767] = 32'hfe5212e3;
        inst_cache[    1768] = 32'h0bc00193;
        inst_cache[    1769] = 32'h00000213;
        inst_cache[    1770] = 32'h00000093;
        inst_cache[    1771] = 32'h00000013;
        inst_cache[    1772] = 32'h00000013;
        inst_cache[    1773] = 32'hfff00113;
        inst_cache[    1774] = 32'h7020c863;
        inst_cache[    1775] = 32'h00120213;
        inst_cache[    1776] = 32'h00200293;
        inst_cache[    1777] = 32'hfe5212e3;
        inst_cache[    1778] = 32'h00100093;
        inst_cache[    1779] = 32'h00104a63;
        inst_cache[    1780] = 32'h00108093;
        inst_cache[    1781] = 32'h00108093;
        inst_cache[    1782] = 32'h00108093;
        inst_cache[    1783] = 32'h00108093;
        inst_cache[    1784] = 32'h00108093;
        inst_cache[    1785] = 32'h00108093;
        inst_cache[    1786] = 32'h00300e93;
        inst_cache[    1787] = 32'h0bd00193;
        inst_cache[    1788] = 32'h6dd09c63;
        inst_cache[    1789] = 32'h0be00193;
        inst_cache[    1790] = 32'h00000093;
        inst_cache[    1791] = 32'h00100113;
        inst_cache[    1792] = 32'h0020e663;
        inst_cache[    1793] = 32'h6c301263;
        inst_cache[    1794] = 32'h00301663;
        inst_cache[    1795] = 32'hfe20eee3;
        inst_cache[    1796] = 32'h6a301c63;
        inst_cache[    1797] = 32'h0bf00193;
        inst_cache[    1798] = 32'hffe00093;
        inst_cache[    1799] = 32'hfff00113;
        inst_cache[    1800] = 32'h0020e663;
        inst_cache[    1801] = 32'h6a301263;
        inst_cache[    1802] = 32'h00301663;
        inst_cache[    1803] = 32'hfe20eee3;
        inst_cache[    1804] = 32'h68301c63;
        inst_cache[    1805] = 32'h0c000193;
        inst_cache[    1806] = 32'h00000093;
        inst_cache[    1807] = 32'hfff00113;
        inst_cache[    1808] = 32'h0020e663;
        inst_cache[    1809] = 32'h68301263;
        inst_cache[    1810] = 32'h00301663;
        inst_cache[    1811] = 32'hfe20eee3;
        inst_cache[    1812] = 32'h66301c63;
        inst_cache[    1813] = 32'h0c100193;
        inst_cache[    1814] = 32'h00100093;
        inst_cache[    1815] = 32'h00000113;
        inst_cache[    1816] = 32'h0020e463;
        inst_cache[    1817] = 32'h00301463;
        inst_cache[    1818] = 32'h66301063;
        inst_cache[    1819] = 32'hfe20eee3;
        inst_cache[    1820] = 32'h0c200193;
        inst_cache[    1821] = 32'hfff00093;
        inst_cache[    1822] = 32'hffe00113;
        inst_cache[    1823] = 32'h0020e463;
        inst_cache[    1824] = 32'h00301463;
        inst_cache[    1825] = 32'h64301263;
        inst_cache[    1826] = 32'hfe20eee3;
        inst_cache[    1827] = 32'h0c300193;
        inst_cache[    1828] = 32'hfff00093;
        inst_cache[    1829] = 32'h00000113;
        inst_cache[    1830] = 32'h0020e463;
        inst_cache[    1831] = 32'h00301463;
        inst_cache[    1832] = 32'h62301463;
        inst_cache[    1833] = 32'hfe20eee3;
        inst_cache[    1834] = 32'h0c400193;
        inst_cache[    1835] = 32'h800000b7;
        inst_cache[    1836] = 32'h80000137;
        inst_cache[    1837] = 32'hfff10113;
        inst_cache[    1838] = 32'h0020e463;
        inst_cache[    1839] = 32'h00301463;
        inst_cache[    1840] = 32'h60301463;
        inst_cache[    1841] = 32'hfe20eee3;
        inst_cache[    1842] = 32'h0c500193;
        inst_cache[    1843] = 32'h00000213;
        inst_cache[    1844] = 32'hf00000b7;
        inst_cache[    1845] = 32'hf0000137;
        inst_cache[    1846] = 32'hfff10113;
        inst_cache[    1847] = 32'h5e20e663;
        inst_cache[    1848] = 32'h00120213;
        inst_cache[    1849] = 32'h00200293;
        inst_cache[    1850] = 32'hfe5214e3;
        inst_cache[    1851] = 32'h0c600193;
        inst_cache[    1852] = 32'h00000213;
        inst_cache[    1853] = 32'hf00000b7;
        inst_cache[    1854] = 32'hf0000137;
        inst_cache[    1855] = 32'hfff10113;
        inst_cache[    1856] = 32'h00000013;
        inst_cache[    1857] = 32'h5c20e263;
        inst_cache[    1858] = 32'h00120213;
        inst_cache[    1859] = 32'h00200293;
        inst_cache[    1860] = 32'hfe5212e3;
        inst_cache[    1861] = 32'h0c700193;
        inst_cache[    1862] = 32'h00000213;
        inst_cache[    1863] = 32'hf00000b7;
        inst_cache[    1864] = 32'hf0000137;
        inst_cache[    1865] = 32'hfff10113;
        inst_cache[    1866] = 32'h00000013;
        inst_cache[    1867] = 32'h00000013;
        inst_cache[    1868] = 32'h5820ec63;
        inst_cache[    1869] = 32'h00120213;
        inst_cache[    1870] = 32'h00200293;
        inst_cache[    1871] = 32'hfe5210e3;
        inst_cache[    1872] = 32'h0c800193;
        inst_cache[    1873] = 32'h00000213;
        inst_cache[    1874] = 32'hf00000b7;
        inst_cache[    1875] = 32'h00000013;
        inst_cache[    1876] = 32'hf0000137;
        inst_cache[    1877] = 32'hfff10113;
        inst_cache[    1878] = 32'h5620e863;
        inst_cache[    1879] = 32'h00120213;
        inst_cache[    1880] = 32'h00200293;
        inst_cache[    1881] = 32'hfe5212e3;
        inst_cache[    1882] = 32'h0c900193;
        inst_cache[    1883] = 32'h00000213;
        inst_cache[    1884] = 32'hf00000b7;
        inst_cache[    1885] = 32'h00000013;
        inst_cache[    1886] = 32'hf0000137;
        inst_cache[    1887] = 32'hfff10113;
        inst_cache[    1888] = 32'h00000013;
        inst_cache[    1889] = 32'h5420e263;
        inst_cache[    1890] = 32'h00120213;
        inst_cache[    1891] = 32'h00200293;
        inst_cache[    1892] = 32'hfe5210e3;
        inst_cache[    1893] = 32'h0ca00193;
        inst_cache[    1894] = 32'h00000213;
        inst_cache[    1895] = 32'hf00000b7;
        inst_cache[    1896] = 32'h00000013;
        inst_cache[    1897] = 32'h00000013;
        inst_cache[    1898] = 32'hf0000137;
        inst_cache[    1899] = 32'hfff10113;
        inst_cache[    1900] = 32'h5020ec63;
        inst_cache[    1901] = 32'h00120213;
        inst_cache[    1902] = 32'h00200293;
        inst_cache[    1903] = 32'hfe5210e3;
        inst_cache[    1904] = 32'h0cb00193;
        inst_cache[    1905] = 32'h00000213;
        inst_cache[    1906] = 32'hf00000b7;
        inst_cache[    1907] = 32'hf0000137;
        inst_cache[    1908] = 32'hfff10113;
        inst_cache[    1909] = 32'h4e20ea63;
        inst_cache[    1910] = 32'h00120213;
        inst_cache[    1911] = 32'h00200293;
        inst_cache[    1912] = 32'hfe5214e3;
        inst_cache[    1913] = 32'h0cc00193;
        inst_cache[    1914] = 32'h00000213;
        inst_cache[    1915] = 32'hf00000b7;
        inst_cache[    1916] = 32'hf0000137;
        inst_cache[    1917] = 32'hfff10113;
        inst_cache[    1918] = 32'h00000013;
        inst_cache[    1919] = 32'h4c20e663;
        inst_cache[    1920] = 32'h00120213;
        inst_cache[    1921] = 32'h00200293;
        inst_cache[    1922] = 32'hfe5212e3;
        inst_cache[    1923] = 32'h0cd00193;
        inst_cache[    1924] = 32'h00000213;
        inst_cache[    1925] = 32'hf00000b7;
        inst_cache[    1926] = 32'hf0000137;
        inst_cache[    1927] = 32'hfff10113;
        inst_cache[    1928] = 32'h00000013;
        inst_cache[    1929] = 32'h00000013;
        inst_cache[    1930] = 32'h4a20e063;
        inst_cache[    1931] = 32'h00120213;
        inst_cache[    1932] = 32'h00200293;
        inst_cache[    1933] = 32'hfe5210e3;
        inst_cache[    1934] = 32'h0ce00193;
        inst_cache[    1935] = 32'h00000213;
        inst_cache[    1936] = 32'hf00000b7;
        inst_cache[    1937] = 32'h00000013;
        inst_cache[    1938] = 32'hf0000137;
        inst_cache[    1939] = 32'hfff10113;
        inst_cache[    1940] = 32'h4620ec63;
        inst_cache[    1941] = 32'h00120213;
        inst_cache[    1942] = 32'h00200293;
        inst_cache[    1943] = 32'hfe5212e3;
        inst_cache[    1944] = 32'h0cf00193;
        inst_cache[    1945] = 32'h00000213;
        inst_cache[    1946] = 32'hf00000b7;
        inst_cache[    1947] = 32'h00000013;
        inst_cache[    1948] = 32'hf0000137;
        inst_cache[    1949] = 32'hfff10113;
        inst_cache[    1950] = 32'h00000013;
        inst_cache[    1951] = 32'h4420e663;
        inst_cache[    1952] = 32'h00120213;
        inst_cache[    1953] = 32'h00200293;
        inst_cache[    1954] = 32'hfe5210e3;
        inst_cache[    1955] = 32'h0d000193;
        inst_cache[    1956] = 32'h00000213;
        inst_cache[    1957] = 32'hf00000b7;
        inst_cache[    1958] = 32'h00000013;
        inst_cache[    1959] = 32'h00000013;
        inst_cache[    1960] = 32'hf0000137;
        inst_cache[    1961] = 32'hfff10113;
        inst_cache[    1962] = 32'h4220e063;
        inst_cache[    1963] = 32'h00120213;
        inst_cache[    1964] = 32'h00200293;
        inst_cache[    1965] = 32'hfe5210e3;
        inst_cache[    1966] = 32'h00100093;
        inst_cache[    1967] = 32'h00106a63;
        inst_cache[    1968] = 32'h00108093;
        inst_cache[    1969] = 32'h00108093;
        inst_cache[    1970] = 32'h00108093;
        inst_cache[    1971] = 32'h00108093;
        inst_cache[    1972] = 32'h00108093;
        inst_cache[    1973] = 32'h00108093;
        inst_cache[    1974] = 32'h00300e93;
        inst_cache[    1975] = 32'h0d100193;
        inst_cache[    1976] = 32'h3fd09463;
        inst_cache[    1977] = 32'h0d200193;
        inst_cache[    1978] = 32'h00000093;
        inst_cache[    1979] = 32'h00100113;
        inst_cache[    1980] = 32'h00209663;
        inst_cache[    1981] = 32'h3c301a63;
        inst_cache[    1982] = 32'h00301663;
        inst_cache[    1983] = 32'hfe209ee3;
        inst_cache[    1984] = 32'h3c301463;
        inst_cache[    1985] = 32'h0d300193;
        inst_cache[    1986] = 32'h00100093;
        inst_cache[    1987] = 32'h00000113;
        inst_cache[    1988] = 32'h00209663;
        inst_cache[    1989] = 32'h3a301a63;
        inst_cache[    1990] = 32'h00301663;
        inst_cache[    1991] = 32'hfe209ee3;
        inst_cache[    1992] = 32'h3a301463;
        inst_cache[    1993] = 32'h0d400193;
        inst_cache[    1994] = 32'hfff00093;
        inst_cache[    1995] = 32'h00100113;
        inst_cache[    1996] = 32'h00209663;
        inst_cache[    1997] = 32'h38301a63;
        inst_cache[    1998] = 32'h00301663;
        inst_cache[    1999] = 32'hfe209ee3;
        inst_cache[    2000] = 32'h38301463;
        inst_cache[    2001] = 32'h0d500193;
        inst_cache[    2002] = 32'h00100093;
        inst_cache[    2003] = 32'hfff00113;
        inst_cache[    2004] = 32'h00209663;
        inst_cache[    2005] = 32'h36301a63;
        inst_cache[    2006] = 32'h00301663;
        inst_cache[    2007] = 32'hfe209ee3;
        inst_cache[    2008] = 32'h36301463;
        inst_cache[    2009] = 32'h0d600193;
        inst_cache[    2010] = 32'h00000093;
        inst_cache[    2011] = 32'h00000113;
        inst_cache[    2012] = 32'h00209463;
        inst_cache[    2013] = 32'h00301463;
        inst_cache[    2014] = 32'h34301863;
        inst_cache[    2015] = 32'hfe209ee3;
        inst_cache[    2016] = 32'h0d700193;
        inst_cache[    2017] = 32'h00100093;
        inst_cache[    2018] = 32'h00100113;
        inst_cache[    2019] = 32'h00209463;
        inst_cache[    2020] = 32'h00301463;
        inst_cache[    2021] = 32'h32301a63;
        inst_cache[    2022] = 32'hfe209ee3;
        inst_cache[    2023] = 32'h0d800193;
        inst_cache[    2024] = 32'hfff00093;
        inst_cache[    2025] = 32'hfff00113;
        inst_cache[    2026] = 32'h00209463;
        inst_cache[    2027] = 32'h00301463;
        inst_cache[    2028] = 32'h30301c63;
        inst_cache[    2029] = 32'hfe209ee3;
        inst_cache[    2030] = 32'h0d900193;
        inst_cache[    2031] = 32'h00000213;
        inst_cache[    2032] = 32'h00000093;
        inst_cache[    2033] = 32'h00000113;
        inst_cache[    2034] = 32'h30209063;
        inst_cache[    2035] = 32'h00120213;
        inst_cache[    2036] = 32'h00200293;
        inst_cache[    2037] = 32'hfe5216e3;
        inst_cache[    2038] = 32'h0da00193;
        inst_cache[    2039] = 32'h00000213;
        inst_cache[    2040] = 32'h00000093;
        inst_cache[    2041] = 32'h00000113;
        inst_cache[    2042] = 32'h00000013;
        inst_cache[    2043] = 32'h2c209e63;
        inst_cache[    2044] = 32'h00120213;
        inst_cache[    2045] = 32'h00200293;
        inst_cache[    2046] = 32'hfe5214e3;
        inst_cache[    2047] = 32'h0db00193;
        inst_cache[    2048] = 32'h00000213;
        inst_cache[    2049] = 32'h00000093;
        inst_cache[    2050] = 32'h00000113;
        inst_cache[    2051] = 32'h00000013;
        inst_cache[    2052] = 32'h00000013;
        inst_cache[    2053] = 32'h2a209a63;
        inst_cache[    2054] = 32'h00120213;
        inst_cache[    2055] = 32'h00200293;
        inst_cache[    2056] = 32'hfe5212e3;
        inst_cache[    2057] = 32'h0dc00193;
        inst_cache[    2058] = 32'h00000213;
        inst_cache[    2059] = 32'h00000093;
        inst_cache[    2060] = 32'h00000013;
        inst_cache[    2061] = 32'h00000113;
        inst_cache[    2062] = 32'h28209863;
        inst_cache[    2063] = 32'h00120213;
        inst_cache[    2064] = 32'h00200293;
        inst_cache[    2065] = 32'hfe5214e3;
        inst_cache[    2066] = 32'h0dd00193;
        inst_cache[    2067] = 32'h00000213;
        inst_cache[    2068] = 32'h00000093;
        inst_cache[    2069] = 32'h00000013;
        inst_cache[    2070] = 32'h00000113;
        inst_cache[    2071] = 32'h00000013;
        inst_cache[    2072] = 32'h26209463;
        inst_cache[    2073] = 32'h00120213;
        inst_cache[    2074] = 32'h00200293;
        inst_cache[    2075] = 32'hfe5212e3;
        inst_cache[    2076] = 32'h0de00193;
        inst_cache[    2077] = 32'h00000213;
        inst_cache[    2078] = 32'h00000093;
        inst_cache[    2079] = 32'h00000013;
        inst_cache[    2080] = 32'h00000013;
        inst_cache[    2081] = 32'h00000113;
        inst_cache[    2082] = 32'h24209063;
        inst_cache[    2083] = 32'h00120213;
        inst_cache[    2084] = 32'h00200293;
        inst_cache[    2085] = 32'hfe5212e3;
        inst_cache[    2086] = 32'h0df00193;
        inst_cache[    2087] = 32'h00000213;
        inst_cache[    2088] = 32'h00000093;
        inst_cache[    2089] = 32'h00000113;
        inst_cache[    2090] = 32'h22209063;
        inst_cache[    2091] = 32'h00120213;
        inst_cache[    2092] = 32'h00200293;
        inst_cache[    2093] = 32'hfe5216e3;
        inst_cache[    2094] = 32'h0e000193;
        inst_cache[    2095] = 32'h00000213;
        inst_cache[    2096] = 32'h00000093;
        inst_cache[    2097] = 32'h00000113;
        inst_cache[    2098] = 32'h00000013;
        inst_cache[    2099] = 32'h1e209e63;
        inst_cache[    2100] = 32'h00120213;
        inst_cache[    2101] = 32'h00200293;
        inst_cache[    2102] = 32'hfe5214e3;
        inst_cache[    2103] = 32'h0e100193;
        inst_cache[    2104] = 32'h00000213;
        inst_cache[    2105] = 32'h00000093;
        inst_cache[    2106] = 32'h00000113;
        inst_cache[    2107] = 32'h00000013;
        inst_cache[    2108] = 32'h00000013;
        inst_cache[    2109] = 32'h1c209a63;
        inst_cache[    2110] = 32'h00120213;
        inst_cache[    2111] = 32'h00200293;
        inst_cache[    2112] = 32'hfe5212e3;
        inst_cache[    2113] = 32'h0e200193;
        inst_cache[    2114] = 32'h00000213;
        inst_cache[    2115] = 32'h00000093;
        inst_cache[    2116] = 32'h00000013;
        inst_cache[    2117] = 32'h00000113;
        inst_cache[    2118] = 32'h1a209863;
        inst_cache[    2119] = 32'h00120213;
        inst_cache[    2120] = 32'h00200293;
        inst_cache[    2121] = 32'hfe5214e3;
        inst_cache[    2122] = 32'h0e300193;
        inst_cache[    2123] = 32'h00000213;
        inst_cache[    2124] = 32'h00000093;
        inst_cache[    2125] = 32'h00000013;
        inst_cache[    2126] = 32'h00000113;
        inst_cache[    2127] = 32'h00000013;
        inst_cache[    2128] = 32'h18209463;
        inst_cache[    2129] = 32'h00120213;
        inst_cache[    2130] = 32'h00200293;
        inst_cache[    2131] = 32'hfe5212e3;
        inst_cache[    2132] = 32'h0e400193;
        inst_cache[    2133] = 32'h00000213;
        inst_cache[    2134] = 32'h00000093;
        inst_cache[    2135] = 32'h00000013;
        inst_cache[    2136] = 32'h00000013;
        inst_cache[    2137] = 32'h00000113;
        inst_cache[    2138] = 32'h16209063;
        inst_cache[    2139] = 32'h00120213;
        inst_cache[    2140] = 32'h00200293;
        inst_cache[    2141] = 32'hfe5212e3;
        inst_cache[    2142] = 32'h00100093;
        inst_cache[    2143] = 32'h00009a63;
        inst_cache[    2144] = 32'h00108093;
        inst_cache[    2145] = 32'h00108093;
        inst_cache[    2146] = 32'h00108093;
        inst_cache[    2147] = 32'h00108093;
        inst_cache[    2148] = 32'h00108093;
        inst_cache[    2149] = 32'h00108093;
        inst_cache[    2150] = 32'h00300e93;
        inst_cache[    2151] = 32'h0e500193;
        inst_cache[    2152] = 32'h13d09463;
        inst_cache[    2153] = 32'h00200193;
        inst_cache[    2154] = 32'h00000093;
        inst_cache[    2155] = 32'h0100026f;
        inst_cache[    2156] = 32'h00000013;
        inst_cache[    2157] = 32'h00000013;
        inst_cache[    2158] = 32'h1100006f;
        inst_cache[    2159] = 32'h00000317;
        inst_cache[    2160] = 32'hff430313;
        inst_cache[    2161] = 32'h10431263;
        inst_cache[    2162] = 32'h00100093;
        inst_cache[    2163] = 32'h0140006f;
        inst_cache[    2164] = 32'h00108093;
        inst_cache[    2165] = 32'h00108093;
        inst_cache[    2166] = 32'h00108093;
        inst_cache[    2167] = 32'h00108093;
        inst_cache[    2168] = 32'h00108093;
        inst_cache[    2169] = 32'h00108093;
        inst_cache[    2170] = 32'h00300e93;
        inst_cache[    2171] = 32'h0e800193;
        inst_cache[    2172] = 32'h0dd09c63;
        inst_cache[    2173] = 32'h00200193;
        inst_cache[    2174] = 32'h00000293;
        inst_cache[    2175] = 32'h00000317;
        inst_cache[    2176] = 32'h01030313;
        inst_cache[    2177] = 32'h000302e7;
        inst_cache[    2178] = 32'h0c00006f;
        inst_cache[    2179] = 32'h00000317;
        inst_cache[    2180] = 32'hffc30313;
        inst_cache[    2181] = 32'h0a629a63;
        inst_cache[    2182] = 32'h0e900193;
        inst_cache[    2183] = 32'h00000213;
        inst_cache[    2184] = 32'h00000317;
        inst_cache[    2185] = 32'h01030313;
        inst_cache[    2186] = 32'h000309e7;
        inst_cache[    2187] = 32'h08301e63;
        inst_cache[    2188] = 32'h00120213;
        inst_cache[    2189] = 32'h00200293;
        inst_cache[    2190] = 32'hfe5214e3;
        inst_cache[    2191] = 32'h0ea00193;
        inst_cache[    2192] = 32'h00000213;
        inst_cache[    2193] = 32'h00000317;
        inst_cache[    2194] = 32'h01430313;
        inst_cache[    2195] = 32'h00000013;
        inst_cache[    2196] = 32'h000309e7;
        inst_cache[    2197] = 32'h06301a63;
        inst_cache[    2198] = 32'h00120213;
        inst_cache[    2199] = 32'h00200293;
        inst_cache[    2200] = 32'hfe5212e3;
        inst_cache[    2201] = 32'h0eb00193;
        inst_cache[    2202] = 32'h00000213;
        inst_cache[    2203] = 32'h00000317;
        inst_cache[    2204] = 32'h01830313;
        inst_cache[    2205] = 32'h00000013;
        inst_cache[    2206] = 32'h00000013;
        inst_cache[    2207] = 32'h000309e7;
        inst_cache[    2208] = 32'h04301463;
        inst_cache[    2209] = 32'h00120213;
        inst_cache[    2210] = 32'h00200293;
        inst_cache[    2211] = 32'hfe5210e3;
        inst_cache[    2212] = 32'h00100293;
        inst_cache[    2213] = 32'h00000317;
        inst_cache[    2214] = 32'h01c30313;
        inst_cache[    2215] = 32'hffc30067;
        inst_cache[    2216] = 32'h00128293;
        inst_cache[    2217] = 32'h00128293;
        inst_cache[    2218] = 32'h00128293;
        inst_cache[    2219] = 32'h00128293;
        inst_cache[    2220] = 32'h00128293;
        inst_cache[    2221] = 32'h00128293;
        inst_cache[    2222] = 32'h00400e93;
        inst_cache[    2223] = 32'h0ec00193;
        inst_cache[    2224] = 32'h01d29463;
        inst_cache[    2225] = 32'h00301463;
        inst_cache[    2226] = 32'h00000a6f;
        inst_cache[    2227] = 32'h00100193;
        inst_cache[    2228] = 32'h00000a6f;
        inst_cache[    2229] = 32'hc0001073;
        inst_cache[    2230] = 32'h00000000;
        inst_cache[    2231] = 32'h00000000;
        inst_cache[    2232] = 32'h00000000;
        inst_cache[    2233] = 32'h00000000;
        inst_cache[    2234] = 32'h00000000;
        inst_cache[    2235] = 32'h00000000;
        inst_cache[    2236] = 32'h00000000;
        inst_cache[    2237] = 32'h00000000;
        inst_cache[    2238] = 32'h00000000;
        inst_cache[    2239] = 32'h00000000;
        inst_cache[    2240] = 32'h00000000;
end
endmodule
